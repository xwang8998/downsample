module rompcm176(
	input clk,//45m
	input reset_n,
	output signed [31:0]addrout
);

wire signed [31:0]addr[0:65535];
reg [7:0]k;
wire lrck;
always @(posedge clk or negedge reset_n)begin
	if(reset_n ==0) 
	k = 0;
	
	else
	k <= k+1;

end
assign lrck = k[7];
reg [15:0]i;
always @(posedge lrck or negedge reset_n)begin
	if(reset_n ==0)begin
		i <= 0;
	//	addrout <= 32'd0;
		end
	
	else begin
		i <= i+1;
	//	addrout <= addr[i];
		end
end

assign addrout = addr[i];
assign addr[0]= 0;
assign addr[1]= 76474970;
assign addr[2]= 152852926;
assign addr[3]= 229036977;
assign addr[4]= 304930476;
assign addr[5]= 380437148;
assign addr[6]= 455461206;
assign addr[7]= 529907477;
assign addr[8]= 603681519;
assign addr[9]= 676689746;
assign addr[10]= 748839539;
assign addr[11]= 820039373;
assign addr[12]= 890198924;
assign addr[13]= 959229189;
assign addr[14]= 1027042599;
assign addr[15]= 1093553126;
assign addr[16]= 1158676398;
assign addr[17]= 1222329801;
assign addr[18]= 1284432584;
assign addr[19]= 1344905966;
assign addr[20]= 1403673233;
assign addr[21]= 1460659832;
assign addr[22]= 1515793473;
assign addr[23]= 1569004214;
assign addr[24]= 1620224553;
assign addr[25]= 1669389513;
assign addr[26]= 1716436725;
assign addr[27]= 1761306505;
assign addr[28]= 1803941934;
assign addr[29]= 1844288924;
assign addr[30]= 1882296293;
assign addr[31]= 1917915825;
assign addr[32]= 1951102334;
assign addr[33]= 1981813720;
assign addr[34]= 2010011024;
assign addr[35]= 2035658475;
assign addr[36]= 2058723538;
assign addr[37]= 2079176953;
assign addr[38]= 2096992772;
assign addr[39]= 2112148396;
assign addr[40]= 2124624598;
assign addr[41]= 2134405552;
assign addr[42]= 2141478848;
assign addr[43]= 2145835515;
assign addr[44]= 2147470025;
assign addr[45]= 2146380306;
assign addr[46]= 2142567738;
assign addr[47]= 2136037160;
assign addr[48]= 2126796855;
assign addr[49]= 2114858546;
assign addr[50]= 2100237377;
assign addr[51]= 2082951896;
assign addr[52]= 2063024031;
assign addr[53]= 2040479063;
assign addr[54]= 2015345591;
assign addr[55]= 1987655498;
assign addr[56]= 1957443913;
assign addr[57]= 1924749160;
assign addr[58]= 1889612716;
assign addr[59]= 1852079154;
assign addr[60]= 1812196087;
assign addr[61]= 1770014111;
assign addr[62]= 1725586737;
assign addr[63]= 1678970324;
assign addr[64]= 1630224009;
assign addr[65]= 1579409630;
assign addr[66]= 1526591649;
assign addr[67]= 1471837070;
assign addr[68]= 1415215352;
assign addr[69]= 1356798326;
assign addr[70]= 1296660098;
assign addr[71]= 1234876957;
assign addr[72]= 1171527280;
assign addr[73]= 1106691431;
assign addr[74]= 1040451659;
assign addr[75]= 972891995;
assign addr[76]= 904098143;
assign addr[77]= 834157373;
assign addr[78]= 763158411;
assign addr[79]= 691191324;
assign addr[80]= 618347408;
assign addr[81]= 544719071;
assign addr[82]= 470399716;
assign addr[83]= 395483624;
assign addr[84]= 320065829;
assign addr[85]= 244242007;
assign addr[86]= 168108346;
assign addr[87]= 91761426;
assign addr[88]= 15298099;
assign addr[89]= -61184634;
assign addr[90]= -137589750;
assign addr[91]= -213820322;
assign addr[92]= -289779648;
assign addr[93]= -365371365;
assign addr[94]= -440499581;
assign addr[95]= -515068990;
assign addr[96]= -588984994;
assign addr[97]= -662153826;
assign addr[98]= -734482665;
assign addr[99]= -805879757;
assign addr[100]= -876254528;
assign addr[101]= -945517704;
assign addr[102]= -1013581418;
assign addr[103]= -1080359326;
assign addr[104]= -1145766716;
assign addr[105]= -1209720613;
assign addr[106]= -1272139887;
assign addr[107]= -1332945355;
assign addr[108]= -1392059879;
assign addr[109]= -1449408469;
assign addr[110]= -1504918373;
assign addr[111]= -1558519173;
assign addr[112]= -1610142873;
assign addr[113]= -1659723983;
assign addr[114]= -1707199606;
assign addr[115]= -1752509516;
assign addr[116]= -1795596234;
assign addr[117]= -1836405100;
assign addr[118]= -1874884346;
assign addr[119]= -1910985158;
assign addr[120]= -1944661739;
assign addr[121]= -1975871368;
assign addr[122]= -2004574453;
assign addr[123]= -2030734582;
assign addr[124]= -2054318569;
assign addr[125]= -2075296495;
assign addr[126]= -2093641749;
assign addr[127]= -2109331059;
assign addr[128]= -2122344521;
assign addr[129]= -2132665626;
assign addr[130]= -2140281282;
assign addr[131]= -2145181827;
assign addr[132]= -2147361045;
assign addr[133]= -2146816171;
assign addr[134]= -2143547897;
assign addr[135]= -2137560369;
assign addr[136]= -2128861181;
assign addr[137]= -2117461370;
assign addr[138]= -2103375398;
assign addr[139]= -2086621133;
assign addr[140]= -2067219829;
assign addr[141]= -2045196100;
assign addr[142]= -2020577882;
assign addr[143]= -1993396407;
assign addr[144]= -1963686155;
assign addr[145]= -1931484818;
assign addr[146]= -1896833245;
assign addr[147]= -1859775393;
assign addr[148]= -1820358275;
assign addr[149]= -1778631892;
assign addr[150]= -1734649179;
assign addr[151]= -1688465931;
assign addr[152]= -1640140734;
assign addr[153]= -1589734894;
assign addr[154]= -1537312353;
assign addr[155]= -1482939614;
assign addr[156]= -1426685652;
assign addr[157]= -1368621831;
assign addr[158]= -1308821808;
assign addr[159]= -1247361445;
assign addr[160]= -1184318708;
assign addr[161]= -1119773573;
assign addr[162]= -1053807919;
assign addr[163]= -986505429;
assign addr[164]= -917951481;
assign addr[165]= -848233042;
assign addr[166]= -777438554;
assign addr[167]= -705657826;
assign addr[168]= -632981917;
assign addr[169]= -559503022;
assign addr[170]= -485314355;
assign addr[171]= -410510029;
assign addr[172]= -335184940;
assign addr[173]= -259434643;
assign addr[174]= -183355234;
assign addr[175]= -107043224;
assign addr[176]= -30595422;
assign addr[177]= 45891193;
assign addr[178]= 122319591;
assign addr[179]= 198592817;
assign addr[180]= 274614114;
assign addr[181]= 350287041;
assign addr[182]= 425515602;
assign addr[183]= 500204365;
assign addr[184]= 574258580;
assign addr[185]= 647584304;
assign addr[186]= 720088517;
assign addr[187]= 791679244;
assign addr[188]= 862265664;
assign addr[189]= 931758235;
assign addr[190]= 1000068799;
assign addr[191]= 1067110699;
assign addr[192]= 1132798888;
assign addr[193]= 1197050035;
assign addr[194]= 1259782632;
assign addr[195]= 1320917099;
assign addr[196]= 1380375881;
assign addr[197]= 1438083551;
assign addr[198]= 1493966902;
assign addr[199]= 1547955041;
assign addr[200]= 1599979481;
assign addr[201]= 1649974225;
assign addr[202]= 1697875851;
assign addr[203]= 1743623590;
assign addr[204]= 1787159411;
assign addr[205]= 1828428082;
assign addr[206]= 1867377253;
assign addr[207]= 1903957513;
assign addr[208]= 1938122457;
assign addr[209]= 1969828744;
assign addr[210]= 1999036154;
assign addr[211]= 2025707632;
assign addr[212]= 2049809346;
assign addr[213]= 2071310720;
assign addr[214]= 2090184478;
assign addr[215]= 2106406677;
assign addr[216]= 2119956737;
assign addr[217]= 2130817471;
assign addr[218]= 2138975100;
assign addr[219]= 2144419275;
assign addr[220]= 2147143090;
assign addr[221]= 2147143090;
assign addr[222]= 2144419275;
assign addr[223]= 2138975100;
assign addr[224]= 2130817471;
assign addr[225]= 2119956737;
assign addr[226]= 2106406677;
assign addr[227]= 2090184478;
assign addr[228]= 2071310720;
assign addr[229]= 2049809346;
assign addr[230]= 2025707632;
assign addr[231]= 1999036154;
assign addr[232]= 1969828744;
assign addr[233]= 1938122457;
assign addr[234]= 1903957513;
assign addr[235]= 1867377253;
assign addr[236]= 1828428082;
assign addr[237]= 1787159411;
assign addr[238]= 1743623590;
assign addr[239]= 1697875851;
assign addr[240]= 1649974225;
assign addr[241]= 1599979481;
assign addr[242]= 1547955041;
assign addr[243]= 1493966902;
assign addr[244]= 1438083551;
assign addr[245]= 1380375881;
assign addr[246]= 1320917099;
assign addr[247]= 1259782632;
assign addr[248]= 1197050035;
assign addr[249]= 1132798888;
assign addr[250]= 1067110699;
assign addr[251]= 1000068799;
assign addr[252]= 931758235;
assign addr[253]= 862265664;
assign addr[254]= 791679244;
assign addr[255]= 720088517;
assign addr[256]= 647584304;
assign addr[257]= 574258580;
assign addr[258]= 500204365;
assign addr[259]= 425515602;
assign addr[260]= 350287041;
assign addr[261]= 274614114;
assign addr[262]= 198592817;
assign addr[263]= 122319591;
assign addr[264]= 45891193;
assign addr[265]= -30595422;
assign addr[266]= -107043224;
assign addr[267]= -183355234;
assign addr[268]= -259434643;
assign addr[269]= -335184940;
assign addr[270]= -410510029;
assign addr[271]= -485314355;
assign addr[272]= -559503022;
assign addr[273]= -632981917;
assign addr[274]= -705657826;
assign addr[275]= -777438554;
assign addr[276]= -848233042;
assign addr[277]= -917951481;
assign addr[278]= -986505429;
assign addr[279]= -1053807919;
assign addr[280]= -1119773573;
assign addr[281]= -1184318708;
assign addr[282]= -1247361445;
assign addr[283]= -1308821808;
assign addr[284]= -1368621831;
assign addr[285]= -1426685652;
assign addr[286]= -1482939614;
assign addr[287]= -1537312353;
assign addr[288]= -1589734894;
assign addr[289]= -1640140734;
assign addr[290]= -1688465931;
assign addr[291]= -1734649179;
assign addr[292]= -1778631892;
assign addr[293]= -1820358275;
assign addr[294]= -1859775393;
assign addr[295]= -1896833245;
assign addr[296]= -1931484818;
assign addr[297]= -1963686155;
assign addr[298]= -1993396407;
assign addr[299]= -2020577882;
assign addr[300]= -2045196100;
assign addr[301]= -2067219829;
assign addr[302]= -2086621133;
assign addr[303]= -2103375398;
assign addr[304]= -2117461370;
assign addr[305]= -2128861181;
assign addr[306]= -2137560369;
assign addr[307]= -2143547897;
assign addr[308]= -2146816171;
assign addr[309]= -2147361045;
assign addr[310]= -2145181827;
assign addr[311]= -2140281282;
assign addr[312]= -2132665626;
assign addr[313]= -2122344521;
assign addr[314]= -2109331059;
assign addr[315]= -2093641749;
assign addr[316]= -2075296495;
assign addr[317]= -2054318569;
assign addr[318]= -2030734582;
assign addr[319]= -2004574453;
assign addr[320]= -1975871368;
assign addr[321]= -1944661739;
assign addr[322]= -1910985158;
assign addr[323]= -1874884346;
assign addr[324]= -1836405100;
assign addr[325]= -1795596234;
assign addr[326]= -1752509516;
assign addr[327]= -1707199606;
assign addr[328]= -1659723983;
assign addr[329]= -1610142873;
assign addr[330]= -1558519173;
assign addr[331]= -1504918373;
assign addr[332]= -1449408469;
assign addr[333]= -1392059879;
assign addr[334]= -1332945355;
assign addr[335]= -1272139887;
assign addr[336]= -1209720613;
assign addr[337]= -1145766716;
assign addr[338]= -1080359326;
assign addr[339]= -1013581418;
assign addr[340]= -945517704;
assign addr[341]= -876254528;
assign addr[342]= -805879757;
assign addr[343]= -734482665;
assign addr[344]= -662153826;
assign addr[345]= -588984994;
assign addr[346]= -515068990;
assign addr[347]= -440499581;
assign addr[348]= -365371365;
assign addr[349]= -289779648;
assign addr[350]= -213820322;
assign addr[351]= -137589750;
assign addr[352]= -61184634;
assign addr[353]= 15298099;
assign addr[354]= 91761426;
assign addr[355]= 168108346;
assign addr[356]= 244242007;
assign addr[357]= 320065829;
assign addr[358]= 395483624;
assign addr[359]= 470399716;
assign addr[360]= 544719071;
assign addr[361]= 618347408;
assign addr[362]= 691191324;
assign addr[363]= 763158411;
assign addr[364]= 834157373;
assign addr[365]= 904098143;
assign addr[366]= 972891995;
assign addr[367]= 1040451659;
assign addr[368]= 1106691431;
assign addr[369]= 1171527280;
assign addr[370]= 1234876957;
assign addr[371]= 1296660098;
assign addr[372]= 1356798326;
assign addr[373]= 1415215352;
assign addr[374]= 1471837070;
assign addr[375]= 1526591649;
assign addr[376]= 1579409630;
assign addr[377]= 1630224009;
assign addr[378]= 1678970324;
assign addr[379]= 1725586737;
assign addr[380]= 1770014111;
assign addr[381]= 1812196087;
assign addr[382]= 1852079154;
assign addr[383]= 1889612716;
assign addr[384]= 1924749160;
assign addr[385]= 1957443913;
assign addr[386]= 1987655498;
assign addr[387]= 2015345591;
assign addr[388]= 2040479063;
assign addr[389]= 2063024031;
assign addr[390]= 2082951896;
assign addr[391]= 2100237377;
assign addr[392]= 2114858546;
assign addr[393]= 2126796855;
assign addr[394]= 2136037160;
assign addr[395]= 2142567738;
assign addr[396]= 2146380306;
assign addr[397]= 2147470025;
assign addr[398]= 2145835515;
assign addr[399]= 2141478848;
assign addr[400]= 2134405552;
assign addr[401]= 2124624598;
assign addr[402]= 2112148396;
assign addr[403]= 2096992772;
assign addr[404]= 2079176953;
assign addr[405]= 2058723538;
assign addr[406]= 2035658475;
assign addr[407]= 2010011024;
assign addr[408]= 1981813720;
assign addr[409]= 1951102334;
assign addr[410]= 1917915825;
assign addr[411]= 1882296293;
assign addr[412]= 1844288924;
assign addr[413]= 1803941934;
assign addr[414]= 1761306505;
assign addr[415]= 1716436725;
assign addr[416]= 1669389513;
assign addr[417]= 1620224553;
assign addr[418]= 1569004214;
assign addr[419]= 1515793473;
assign addr[420]= 1460659832;
assign addr[421]= 1403673233;
assign addr[422]= 1344905966;
assign addr[423]= 1284432584;
assign addr[424]= 1222329801;
assign addr[425]= 1158676398;
assign addr[426]= 1093553126;
assign addr[427]= 1027042599;
assign addr[428]= 959229189;
assign addr[429]= 890198924;
assign addr[430]= 820039373;
assign addr[431]= 748839539;
assign addr[432]= 676689746;
assign addr[433]= 603681519;
assign addr[434]= 529907477;
assign addr[435]= 455461206;
assign addr[436]= 380437148;
assign addr[437]= 304930476;
assign addr[438]= 229036977;
assign addr[439]= 152852926;
assign addr[440]= 76474970;
assign addr[441]= 0;
assign addr[442]= -76474970;
assign addr[443]= -152852926;
assign addr[444]= -229036977;
assign addr[445]= -304930476;
assign addr[446]= -380437148;
assign addr[447]= -455461206;
assign addr[448]= -529907477;
assign addr[449]= -603681519;
assign addr[450]= -676689746;
assign addr[451]= -748839539;
assign addr[452]= -820039373;
assign addr[453]= -890198924;
assign addr[454]= -959229189;
assign addr[455]= -1027042599;
assign addr[456]= -1093553126;
assign addr[457]= -1158676398;
assign addr[458]= -1222329801;
assign addr[459]= -1284432584;
assign addr[460]= -1344905966;
assign addr[461]= -1403673233;
assign addr[462]= -1460659832;
assign addr[463]= -1515793473;
assign addr[464]= -1569004214;
assign addr[465]= -1620224553;
assign addr[466]= -1669389513;
assign addr[467]= -1716436725;
assign addr[468]= -1761306505;
assign addr[469]= -1803941934;
assign addr[470]= -1844288924;
assign addr[471]= -1882296293;
assign addr[472]= -1917915825;
assign addr[473]= -1951102334;
assign addr[474]= -1981813720;
assign addr[475]= -2010011024;
assign addr[476]= -2035658475;
assign addr[477]= -2058723538;
assign addr[478]= -2079176953;
assign addr[479]= -2096992772;
assign addr[480]= -2112148396;
assign addr[481]= -2124624598;
assign addr[482]= -2134405552;
assign addr[483]= -2141478848;
assign addr[484]= -2145835515;
assign addr[485]= -2147470025;
assign addr[486]= -2146380306;
assign addr[487]= -2142567738;
assign addr[488]= -2136037160;
assign addr[489]= -2126796855;
assign addr[490]= -2114858546;
assign addr[491]= -2100237377;
assign addr[492]= -2082951896;
assign addr[493]= -2063024031;
assign addr[494]= -2040479063;
assign addr[495]= -2015345591;
assign addr[496]= -1987655498;
assign addr[497]= -1957443913;
assign addr[498]= -1924749160;
assign addr[499]= -1889612716;
assign addr[500]= -1852079154;
assign addr[501]= -1812196087;
assign addr[502]= -1770014111;
assign addr[503]= -1725586737;
assign addr[504]= -1678970324;
assign addr[505]= -1630224009;
assign addr[506]= -1579409630;
assign addr[507]= -1526591649;
assign addr[508]= -1471837070;
assign addr[509]= -1415215352;
assign addr[510]= -1356798326;
assign addr[511]= -1296660098;
assign addr[512]= -1234876957;
assign addr[513]= -1171527280;
assign addr[514]= -1106691431;
assign addr[515]= -1040451659;
assign addr[516]= -972891995;
assign addr[517]= -904098143;
assign addr[518]= -834157373;
assign addr[519]= -763158411;
assign addr[520]= -691191324;
assign addr[521]= -618347408;
assign addr[522]= -544719071;
assign addr[523]= -470399716;
assign addr[524]= -395483624;
assign addr[525]= -320065829;
assign addr[526]= -244242007;
assign addr[527]= -168108346;
assign addr[528]= -91761426;
assign addr[529]= -15298099;
assign addr[530]= 61184634;
assign addr[531]= 137589750;
assign addr[532]= 213820322;
assign addr[533]= 289779648;
assign addr[534]= 365371365;
assign addr[535]= 440499581;
assign addr[536]= 515068990;
assign addr[537]= 588984994;
assign addr[538]= 662153826;
assign addr[539]= 734482665;
assign addr[540]= 805879757;
assign addr[541]= 876254528;
assign addr[542]= 945517704;
assign addr[543]= 1013581418;
assign addr[544]= 1080359326;
assign addr[545]= 1145766716;
assign addr[546]= 1209720613;
assign addr[547]= 1272139887;
assign addr[548]= 1332945355;
assign addr[549]= 1392059879;
assign addr[550]= 1449408469;
assign addr[551]= 1504918373;
assign addr[552]= 1558519173;
assign addr[553]= 1610142873;
assign addr[554]= 1659723983;
assign addr[555]= 1707199606;
assign addr[556]= 1752509516;
assign addr[557]= 1795596234;
assign addr[558]= 1836405100;
assign addr[559]= 1874884346;
assign addr[560]= 1910985158;
assign addr[561]= 1944661739;
assign addr[562]= 1975871368;
assign addr[563]= 2004574453;
assign addr[564]= 2030734582;
assign addr[565]= 2054318569;
assign addr[566]= 2075296495;
assign addr[567]= 2093641749;
assign addr[568]= 2109331059;
assign addr[569]= 2122344521;
assign addr[570]= 2132665626;
assign addr[571]= 2140281282;
assign addr[572]= 2145181827;
assign addr[573]= 2147361045;
assign addr[574]= 2146816171;
assign addr[575]= 2143547897;
assign addr[576]= 2137560369;
assign addr[577]= 2128861181;
assign addr[578]= 2117461370;
assign addr[579]= 2103375398;
assign addr[580]= 2086621133;
assign addr[581]= 2067219829;
assign addr[582]= 2045196100;
assign addr[583]= 2020577882;
assign addr[584]= 1993396407;
assign addr[585]= 1963686155;
assign addr[586]= 1931484818;
assign addr[587]= 1896833245;
assign addr[588]= 1859775393;
assign addr[589]= 1820358275;
assign addr[590]= 1778631892;
assign addr[591]= 1734649179;
assign addr[592]= 1688465931;
assign addr[593]= 1640140734;
assign addr[594]= 1589734894;
assign addr[595]= 1537312353;
assign addr[596]= 1482939614;
assign addr[597]= 1426685652;
assign addr[598]= 1368621831;
assign addr[599]= 1308821808;
assign addr[600]= 1247361445;
assign addr[601]= 1184318708;
assign addr[602]= 1119773573;
assign addr[603]= 1053807919;
assign addr[604]= 986505429;
assign addr[605]= 917951481;
assign addr[606]= 848233042;
assign addr[607]= 777438554;
assign addr[608]= 705657826;
assign addr[609]= 632981917;
assign addr[610]= 559503022;
assign addr[611]= 485314355;
assign addr[612]= 410510029;
assign addr[613]= 335184940;
assign addr[614]= 259434643;
assign addr[615]= 183355234;
assign addr[616]= 107043224;
assign addr[617]= 30595422;
assign addr[618]= -45891193;
assign addr[619]= -122319591;
assign addr[620]= -198592817;
assign addr[621]= -274614114;
assign addr[622]= -350287041;
assign addr[623]= -425515602;
assign addr[624]= -500204365;
assign addr[625]= -574258580;
assign addr[626]= -647584304;
assign addr[627]= -720088517;
assign addr[628]= -791679244;
assign addr[629]= -862265664;
assign addr[630]= -931758235;
assign addr[631]= -1000068799;
assign addr[632]= -1067110699;
assign addr[633]= -1132798888;
assign addr[634]= -1197050035;
assign addr[635]= -1259782632;
assign addr[636]= -1320917099;
assign addr[637]= -1380375881;
assign addr[638]= -1438083551;
assign addr[639]= -1493966902;
assign addr[640]= -1547955041;
assign addr[641]= -1599979481;
assign addr[642]= -1649974225;
assign addr[643]= -1697875851;
assign addr[644]= -1743623590;
assign addr[645]= -1787159411;
assign addr[646]= -1828428082;
assign addr[647]= -1867377253;
assign addr[648]= -1903957513;
assign addr[649]= -1938122457;
assign addr[650]= -1969828744;
assign addr[651]= -1999036154;
assign addr[652]= -2025707632;
assign addr[653]= -2049809346;
assign addr[654]= -2071310720;
assign addr[655]= -2090184478;
assign addr[656]= -2106406677;
assign addr[657]= -2119956737;
assign addr[658]= -2130817471;
assign addr[659]= -2138975100;
assign addr[660]= -2144419275;
assign addr[661]= -2147143090;
assign addr[662]= -2147143090;
assign addr[663]= -2144419275;
assign addr[664]= -2138975100;
assign addr[665]= -2130817471;
assign addr[666]= -2119956737;
assign addr[667]= -2106406677;
assign addr[668]= -2090184478;
assign addr[669]= -2071310720;
assign addr[670]= -2049809346;
assign addr[671]= -2025707632;
assign addr[672]= -1999036154;
assign addr[673]= -1969828744;
assign addr[674]= -1938122457;
assign addr[675]= -1903957513;
assign addr[676]= -1867377253;
assign addr[677]= -1828428082;
assign addr[678]= -1787159411;
assign addr[679]= -1743623590;
assign addr[680]= -1697875851;
assign addr[681]= -1649974225;
assign addr[682]= -1599979481;
assign addr[683]= -1547955041;
assign addr[684]= -1493966902;
assign addr[685]= -1438083551;
assign addr[686]= -1380375881;
assign addr[687]= -1320917099;
assign addr[688]= -1259782632;
assign addr[689]= -1197050035;
assign addr[690]= -1132798888;
assign addr[691]= -1067110699;
assign addr[692]= -1000068799;
assign addr[693]= -931758235;
assign addr[694]= -862265664;
assign addr[695]= -791679244;
assign addr[696]= -720088517;
assign addr[697]= -647584304;
assign addr[698]= -574258580;
assign addr[699]= -500204365;
assign addr[700]= -425515602;
assign addr[701]= -350287041;
assign addr[702]= -274614114;
assign addr[703]= -198592817;
assign addr[704]= -122319591;
assign addr[705]= -45891193;
assign addr[706]= 30595422;
assign addr[707]= 107043224;
assign addr[708]= 183355234;
assign addr[709]= 259434643;
assign addr[710]= 335184940;
assign addr[711]= 410510029;
assign addr[712]= 485314355;
assign addr[713]= 559503022;
assign addr[714]= 632981917;
assign addr[715]= 705657826;
assign addr[716]= 777438554;
assign addr[717]= 848233042;
assign addr[718]= 917951481;
assign addr[719]= 986505429;
assign addr[720]= 1053807919;
assign addr[721]= 1119773573;
assign addr[722]= 1184318708;
assign addr[723]= 1247361445;
assign addr[724]= 1308821808;
assign addr[725]= 1368621831;
assign addr[726]= 1426685652;
assign addr[727]= 1482939614;
assign addr[728]= 1537312353;
assign addr[729]= 1589734894;
assign addr[730]= 1640140734;
assign addr[731]= 1688465931;
assign addr[732]= 1734649179;
assign addr[733]= 1778631892;
assign addr[734]= 1820358275;
assign addr[735]= 1859775393;
assign addr[736]= 1896833245;
assign addr[737]= 1931484818;
assign addr[738]= 1963686155;
assign addr[739]= 1993396407;
assign addr[740]= 2020577882;
assign addr[741]= 2045196100;
assign addr[742]= 2067219829;
assign addr[743]= 2086621133;
assign addr[744]= 2103375398;
assign addr[745]= 2117461370;
assign addr[746]= 2128861181;
assign addr[747]= 2137560369;
assign addr[748]= 2143547897;
assign addr[749]= 2146816171;
assign addr[750]= 2147361045;
assign addr[751]= 2145181827;
assign addr[752]= 2140281282;
assign addr[753]= 2132665626;
assign addr[754]= 2122344521;
assign addr[755]= 2109331059;
assign addr[756]= 2093641749;
assign addr[757]= 2075296495;
assign addr[758]= 2054318569;
assign addr[759]= 2030734582;
assign addr[760]= 2004574453;
assign addr[761]= 1975871368;
assign addr[762]= 1944661739;
assign addr[763]= 1910985158;
assign addr[764]= 1874884346;
assign addr[765]= 1836405100;
assign addr[766]= 1795596234;
assign addr[767]= 1752509516;
assign addr[768]= 1707199606;
assign addr[769]= 1659723983;
assign addr[770]= 1610142873;
assign addr[771]= 1558519173;
assign addr[772]= 1504918373;
assign addr[773]= 1449408469;
assign addr[774]= 1392059879;
assign addr[775]= 1332945355;
assign addr[776]= 1272139887;
assign addr[777]= 1209720613;
assign addr[778]= 1145766716;
assign addr[779]= 1080359326;
assign addr[780]= 1013581418;
assign addr[781]= 945517704;
assign addr[782]= 876254528;
assign addr[783]= 805879757;
assign addr[784]= 734482665;
assign addr[785]= 662153826;
assign addr[786]= 588984994;
assign addr[787]= 515068990;
assign addr[788]= 440499581;
assign addr[789]= 365371365;
assign addr[790]= 289779648;
assign addr[791]= 213820322;
assign addr[792]= 137589750;
assign addr[793]= 61184634;
assign addr[794]= -15298099;
assign addr[795]= -91761426;
assign addr[796]= -168108346;
assign addr[797]= -244242007;
assign addr[798]= -320065829;
assign addr[799]= -395483624;
assign addr[800]= -470399716;
assign addr[801]= -544719071;
assign addr[802]= -618347408;
assign addr[803]= -691191324;
assign addr[804]= -763158411;
assign addr[805]= -834157373;
assign addr[806]= -904098143;
assign addr[807]= -972891995;
assign addr[808]= -1040451659;
assign addr[809]= -1106691431;
assign addr[810]= -1171527280;
assign addr[811]= -1234876957;
assign addr[812]= -1296660098;
assign addr[813]= -1356798326;
assign addr[814]= -1415215352;
assign addr[815]= -1471837070;
assign addr[816]= -1526591649;
assign addr[817]= -1579409630;
assign addr[818]= -1630224009;
assign addr[819]= -1678970324;
assign addr[820]= -1725586737;
assign addr[821]= -1770014111;
assign addr[822]= -1812196087;
assign addr[823]= -1852079154;
assign addr[824]= -1889612716;
assign addr[825]= -1924749160;
assign addr[826]= -1957443913;
assign addr[827]= -1987655498;
assign addr[828]= -2015345591;
assign addr[829]= -2040479063;
assign addr[830]= -2063024031;
assign addr[831]= -2082951896;
assign addr[832]= -2100237377;
assign addr[833]= -2114858546;
assign addr[834]= -2126796855;
assign addr[835]= -2136037160;
assign addr[836]= -2142567738;
assign addr[837]= -2146380306;
assign addr[838]= -2147470025;
assign addr[839]= -2145835515;
assign addr[840]= -2141478848;
assign addr[841]= -2134405552;
assign addr[842]= -2124624598;
assign addr[843]= -2112148396;
assign addr[844]= -2096992772;
assign addr[845]= -2079176953;
assign addr[846]= -2058723538;
assign addr[847]= -2035658475;
assign addr[848]= -2010011024;
assign addr[849]= -1981813720;
assign addr[850]= -1951102334;
assign addr[851]= -1917915825;
assign addr[852]= -1882296293;
assign addr[853]= -1844288924;
assign addr[854]= -1803941934;
assign addr[855]= -1761306505;
assign addr[856]= -1716436725;
assign addr[857]= -1669389513;
assign addr[858]= -1620224553;
assign addr[859]= -1569004214;
assign addr[860]= -1515793473;
assign addr[861]= -1460659832;
assign addr[862]= -1403673233;
assign addr[863]= -1344905966;
assign addr[864]= -1284432584;
assign addr[865]= -1222329801;
assign addr[866]= -1158676398;
assign addr[867]= -1093553126;
assign addr[868]= -1027042599;
assign addr[869]= -959229189;
assign addr[870]= -890198924;
assign addr[871]= -820039373;
assign addr[872]= -748839539;
assign addr[873]= -676689746;
assign addr[874]= -603681519;
assign addr[875]= -529907477;
assign addr[876]= -455461206;
assign addr[877]= -380437148;
assign addr[878]= -304930476;
assign addr[879]= -229036977;
assign addr[880]= -152852926;
assign addr[881]= -76474970;
assign addr[882]= 0;
assign addr[883]= 76474970;
assign addr[884]= 152852926;
assign addr[885]= 229036977;
assign addr[886]= 304930476;
assign addr[887]= 380437148;
assign addr[888]= 455461206;
assign addr[889]= 529907477;
assign addr[890]= 603681519;
assign addr[891]= 676689746;
assign addr[892]= 748839539;
assign addr[893]= 820039373;
assign addr[894]= 890198924;
assign addr[895]= 959229189;
assign addr[896]= 1027042599;
assign addr[897]= 1093553126;
assign addr[898]= 1158676398;
assign addr[899]= 1222329801;
assign addr[900]= 1284432584;
assign addr[901]= 1344905966;
assign addr[902]= 1403673233;
assign addr[903]= 1460659832;
assign addr[904]= 1515793473;
assign addr[905]= 1569004214;
assign addr[906]= 1620224553;
assign addr[907]= 1669389513;
assign addr[908]= 1716436725;
assign addr[909]= 1761306505;
assign addr[910]= 1803941934;
assign addr[911]= 1844288924;
assign addr[912]= 1882296293;
assign addr[913]= 1917915825;
assign addr[914]= 1951102334;
assign addr[915]= 1981813720;
assign addr[916]= 2010011024;
assign addr[917]= 2035658475;
assign addr[918]= 2058723538;
assign addr[919]= 2079176953;
assign addr[920]= 2096992772;
assign addr[921]= 2112148396;
assign addr[922]= 2124624598;
assign addr[923]= 2134405552;
assign addr[924]= 2141478848;
assign addr[925]= 2145835515;
assign addr[926]= 2147470025;
assign addr[927]= 2146380306;
assign addr[928]= 2142567738;
assign addr[929]= 2136037160;
assign addr[930]= 2126796855;
assign addr[931]= 2114858546;
assign addr[932]= 2100237377;
assign addr[933]= 2082951896;
assign addr[934]= 2063024031;
assign addr[935]= 2040479063;
assign addr[936]= 2015345591;
assign addr[937]= 1987655498;
assign addr[938]= 1957443913;
assign addr[939]= 1924749160;
assign addr[940]= 1889612716;
assign addr[941]= 1852079154;
assign addr[942]= 1812196087;
assign addr[943]= 1770014111;
assign addr[944]= 1725586737;
assign addr[945]= 1678970324;
assign addr[946]= 1630224009;
assign addr[947]= 1579409630;
assign addr[948]= 1526591649;
assign addr[949]= 1471837070;
assign addr[950]= 1415215352;
assign addr[951]= 1356798326;
assign addr[952]= 1296660098;
assign addr[953]= 1234876957;
assign addr[954]= 1171527280;
assign addr[955]= 1106691431;
assign addr[956]= 1040451659;
assign addr[957]= 972891995;
assign addr[958]= 904098143;
assign addr[959]= 834157373;
assign addr[960]= 763158411;
assign addr[961]= 691191324;
assign addr[962]= 618347408;
assign addr[963]= 544719071;
assign addr[964]= 470399716;
assign addr[965]= 395483624;
assign addr[966]= 320065829;
assign addr[967]= 244242007;
assign addr[968]= 168108346;
assign addr[969]= 91761426;
assign addr[970]= 15298099;
assign addr[971]= -61184634;
assign addr[972]= -137589750;
assign addr[973]= -213820322;
assign addr[974]= -289779648;
assign addr[975]= -365371365;
assign addr[976]= -440499581;
assign addr[977]= -515068990;
assign addr[978]= -588984994;
assign addr[979]= -662153826;
assign addr[980]= -734482665;
assign addr[981]= -805879757;
assign addr[982]= -876254528;
assign addr[983]= -945517704;
assign addr[984]= -1013581418;
assign addr[985]= -1080359326;
assign addr[986]= -1145766716;
assign addr[987]= -1209720613;
assign addr[988]= -1272139887;
assign addr[989]= -1332945355;
assign addr[990]= -1392059879;
assign addr[991]= -1449408469;
assign addr[992]= -1504918373;
assign addr[993]= -1558519173;
assign addr[994]= -1610142873;
assign addr[995]= -1659723983;
assign addr[996]= -1707199606;
assign addr[997]= -1752509516;
assign addr[998]= -1795596234;
assign addr[999]= -1836405100;
assign addr[1000]= -1874884346;
assign addr[1001]= -1910985158;
assign addr[1002]= -1944661739;
assign addr[1003]= -1975871368;
assign addr[1004]= -2004574453;
assign addr[1005]= -2030734582;
assign addr[1006]= -2054318569;
assign addr[1007]= -2075296495;
assign addr[1008]= -2093641749;
assign addr[1009]= -2109331059;
assign addr[1010]= -2122344521;
assign addr[1011]= -2132665626;
assign addr[1012]= -2140281282;
assign addr[1013]= -2145181827;
assign addr[1014]= -2147361045;
assign addr[1015]= -2146816171;
assign addr[1016]= -2143547897;
assign addr[1017]= -2137560369;
assign addr[1018]= -2128861181;
assign addr[1019]= -2117461370;
assign addr[1020]= -2103375398;
assign addr[1021]= -2086621133;
assign addr[1022]= -2067219829;
assign addr[1023]= -2045196100;
assign addr[1024]= -2020577882;
assign addr[1025]= -1993396407;
assign addr[1026]= -1963686155;
assign addr[1027]= -1931484818;
assign addr[1028]= -1896833245;
assign addr[1029]= -1859775393;
assign addr[1030]= -1820358275;
assign addr[1031]= -1778631892;
assign addr[1032]= -1734649179;
assign addr[1033]= -1688465931;
assign addr[1034]= -1640140734;
assign addr[1035]= -1589734894;
assign addr[1036]= -1537312353;
assign addr[1037]= -1482939614;
assign addr[1038]= -1426685652;
assign addr[1039]= -1368621831;
assign addr[1040]= -1308821808;
assign addr[1041]= -1247361445;
assign addr[1042]= -1184318708;
assign addr[1043]= -1119773573;
assign addr[1044]= -1053807919;
assign addr[1045]= -986505429;
assign addr[1046]= -917951481;
assign addr[1047]= -848233042;
assign addr[1048]= -777438554;
assign addr[1049]= -705657826;
assign addr[1050]= -632981917;
assign addr[1051]= -559503022;
assign addr[1052]= -485314355;
assign addr[1053]= -410510029;
assign addr[1054]= -335184940;
assign addr[1055]= -259434643;
assign addr[1056]= -183355234;
assign addr[1057]= -107043224;
assign addr[1058]= -30595422;
assign addr[1059]= 45891193;
assign addr[1060]= 122319591;
assign addr[1061]= 198592817;
assign addr[1062]= 274614114;
assign addr[1063]= 350287041;
assign addr[1064]= 425515602;
assign addr[1065]= 500204365;
assign addr[1066]= 574258580;
assign addr[1067]= 647584304;
assign addr[1068]= 720088517;
assign addr[1069]= 791679244;
assign addr[1070]= 862265664;
assign addr[1071]= 931758235;
assign addr[1072]= 1000068799;
assign addr[1073]= 1067110699;
assign addr[1074]= 1132798888;
assign addr[1075]= 1197050035;
assign addr[1076]= 1259782632;
assign addr[1077]= 1320917099;
assign addr[1078]= 1380375881;
assign addr[1079]= 1438083551;
assign addr[1080]= 1493966902;
assign addr[1081]= 1547955041;
assign addr[1082]= 1599979481;
assign addr[1083]= 1649974225;
assign addr[1084]= 1697875851;
assign addr[1085]= 1743623590;
assign addr[1086]= 1787159411;
assign addr[1087]= 1828428082;
assign addr[1088]= 1867377253;
assign addr[1089]= 1903957513;
assign addr[1090]= 1938122457;
assign addr[1091]= 1969828744;
assign addr[1092]= 1999036154;
assign addr[1093]= 2025707632;
assign addr[1094]= 2049809346;
assign addr[1095]= 2071310720;
assign addr[1096]= 2090184478;
assign addr[1097]= 2106406677;
assign addr[1098]= 2119956737;
assign addr[1099]= 2130817471;
assign addr[1100]= 2138975100;
assign addr[1101]= 2144419275;
assign addr[1102]= 2147143090;
assign addr[1103]= 2147143090;
assign addr[1104]= 2144419275;
assign addr[1105]= 2138975100;
assign addr[1106]= 2130817471;
assign addr[1107]= 2119956737;
assign addr[1108]= 2106406677;
assign addr[1109]= 2090184478;
assign addr[1110]= 2071310720;
assign addr[1111]= 2049809346;
assign addr[1112]= 2025707632;
assign addr[1113]= 1999036154;
assign addr[1114]= 1969828744;
assign addr[1115]= 1938122457;
assign addr[1116]= 1903957513;
assign addr[1117]= 1867377253;
assign addr[1118]= 1828428082;
assign addr[1119]= 1787159411;
assign addr[1120]= 1743623590;
assign addr[1121]= 1697875851;
assign addr[1122]= 1649974225;
assign addr[1123]= 1599979481;
assign addr[1124]= 1547955041;
assign addr[1125]= 1493966902;
assign addr[1126]= 1438083551;
assign addr[1127]= 1380375881;
assign addr[1128]= 1320917099;
assign addr[1129]= 1259782632;
assign addr[1130]= 1197050035;
assign addr[1131]= 1132798888;
assign addr[1132]= 1067110699;
assign addr[1133]= 1000068799;
assign addr[1134]= 931758235;
assign addr[1135]= 862265664;
assign addr[1136]= 791679244;
assign addr[1137]= 720088517;
assign addr[1138]= 647584304;
assign addr[1139]= 574258580;
assign addr[1140]= 500204365;
assign addr[1141]= 425515602;
assign addr[1142]= 350287041;
assign addr[1143]= 274614114;
assign addr[1144]= 198592817;
assign addr[1145]= 122319591;
assign addr[1146]= 45891193;
assign addr[1147]= -30595422;
assign addr[1148]= -107043224;
assign addr[1149]= -183355234;
assign addr[1150]= -259434643;
assign addr[1151]= -335184940;
assign addr[1152]= -410510029;
assign addr[1153]= -485314355;
assign addr[1154]= -559503022;
assign addr[1155]= -632981917;
assign addr[1156]= -705657826;
assign addr[1157]= -777438554;
assign addr[1158]= -848233042;
assign addr[1159]= -917951481;
assign addr[1160]= -986505429;
assign addr[1161]= -1053807919;
assign addr[1162]= -1119773573;
assign addr[1163]= -1184318708;
assign addr[1164]= -1247361445;
assign addr[1165]= -1308821808;
assign addr[1166]= -1368621831;
assign addr[1167]= -1426685652;
assign addr[1168]= -1482939614;
assign addr[1169]= -1537312353;
assign addr[1170]= -1589734894;
assign addr[1171]= -1640140734;
assign addr[1172]= -1688465931;
assign addr[1173]= -1734649179;
assign addr[1174]= -1778631892;
assign addr[1175]= -1820358275;
assign addr[1176]= -1859775393;
assign addr[1177]= -1896833245;
assign addr[1178]= -1931484818;
assign addr[1179]= -1963686155;
assign addr[1180]= -1993396407;
assign addr[1181]= -2020577882;
assign addr[1182]= -2045196100;
assign addr[1183]= -2067219829;
assign addr[1184]= -2086621133;
assign addr[1185]= -2103375398;
assign addr[1186]= -2117461370;
assign addr[1187]= -2128861181;
assign addr[1188]= -2137560369;
assign addr[1189]= -2143547897;
assign addr[1190]= -2146816171;
assign addr[1191]= -2147361045;
assign addr[1192]= -2145181827;
assign addr[1193]= -2140281282;
assign addr[1194]= -2132665626;
assign addr[1195]= -2122344521;
assign addr[1196]= -2109331059;
assign addr[1197]= -2093641749;
assign addr[1198]= -2075296495;
assign addr[1199]= -2054318569;
assign addr[1200]= -2030734582;
assign addr[1201]= -2004574453;
assign addr[1202]= -1975871368;
assign addr[1203]= -1944661739;
assign addr[1204]= -1910985158;
assign addr[1205]= -1874884346;
assign addr[1206]= -1836405100;
assign addr[1207]= -1795596234;
assign addr[1208]= -1752509516;
assign addr[1209]= -1707199606;
assign addr[1210]= -1659723983;
assign addr[1211]= -1610142873;
assign addr[1212]= -1558519173;
assign addr[1213]= -1504918373;
assign addr[1214]= -1449408469;
assign addr[1215]= -1392059879;
assign addr[1216]= -1332945355;
assign addr[1217]= -1272139887;
assign addr[1218]= -1209720613;
assign addr[1219]= -1145766716;
assign addr[1220]= -1080359326;
assign addr[1221]= -1013581418;
assign addr[1222]= -945517704;
assign addr[1223]= -876254528;
assign addr[1224]= -805879757;
assign addr[1225]= -734482665;
assign addr[1226]= -662153826;
assign addr[1227]= -588984994;
assign addr[1228]= -515068990;
assign addr[1229]= -440499581;
assign addr[1230]= -365371365;
assign addr[1231]= -289779648;
assign addr[1232]= -213820322;
assign addr[1233]= -137589750;
assign addr[1234]= -61184634;
assign addr[1235]= 15298099;
assign addr[1236]= 91761426;
assign addr[1237]= 168108346;
assign addr[1238]= 244242007;
assign addr[1239]= 320065829;
assign addr[1240]= 395483624;
assign addr[1241]= 470399716;
assign addr[1242]= 544719071;
assign addr[1243]= 618347408;
assign addr[1244]= 691191324;
assign addr[1245]= 763158411;
assign addr[1246]= 834157373;
assign addr[1247]= 904098143;
assign addr[1248]= 972891995;
assign addr[1249]= 1040451659;
assign addr[1250]= 1106691431;
assign addr[1251]= 1171527280;
assign addr[1252]= 1234876957;
assign addr[1253]= 1296660098;
assign addr[1254]= 1356798326;
assign addr[1255]= 1415215352;
assign addr[1256]= 1471837070;
assign addr[1257]= 1526591649;
assign addr[1258]= 1579409630;
assign addr[1259]= 1630224009;
assign addr[1260]= 1678970324;
assign addr[1261]= 1725586737;
assign addr[1262]= 1770014111;
assign addr[1263]= 1812196087;
assign addr[1264]= 1852079154;
assign addr[1265]= 1889612716;
assign addr[1266]= 1924749160;
assign addr[1267]= 1957443913;
assign addr[1268]= 1987655498;
assign addr[1269]= 2015345591;
assign addr[1270]= 2040479063;
assign addr[1271]= 2063024031;
assign addr[1272]= 2082951896;
assign addr[1273]= 2100237377;
assign addr[1274]= 2114858546;
assign addr[1275]= 2126796855;
assign addr[1276]= 2136037160;
assign addr[1277]= 2142567738;
assign addr[1278]= 2146380306;
assign addr[1279]= 2147470025;
assign addr[1280]= 2145835515;
assign addr[1281]= 2141478848;
assign addr[1282]= 2134405552;
assign addr[1283]= 2124624598;
assign addr[1284]= 2112148396;
assign addr[1285]= 2096992772;
assign addr[1286]= 2079176953;
assign addr[1287]= 2058723538;
assign addr[1288]= 2035658475;
assign addr[1289]= 2010011024;
assign addr[1290]= 1981813720;
assign addr[1291]= 1951102334;
assign addr[1292]= 1917915825;
assign addr[1293]= 1882296293;
assign addr[1294]= 1844288924;
assign addr[1295]= 1803941934;
assign addr[1296]= 1761306505;
assign addr[1297]= 1716436725;
assign addr[1298]= 1669389513;
assign addr[1299]= 1620224553;
assign addr[1300]= 1569004214;
assign addr[1301]= 1515793473;
assign addr[1302]= 1460659832;
assign addr[1303]= 1403673233;
assign addr[1304]= 1344905966;
assign addr[1305]= 1284432584;
assign addr[1306]= 1222329801;
assign addr[1307]= 1158676398;
assign addr[1308]= 1093553126;
assign addr[1309]= 1027042599;
assign addr[1310]= 959229189;
assign addr[1311]= 890198924;
assign addr[1312]= 820039373;
assign addr[1313]= 748839539;
assign addr[1314]= 676689746;
assign addr[1315]= 603681519;
assign addr[1316]= 529907477;
assign addr[1317]= 455461206;
assign addr[1318]= 380437148;
assign addr[1319]= 304930476;
assign addr[1320]= 229036977;
assign addr[1321]= 152852926;
assign addr[1322]= 76474970;
assign addr[1323]= 0;
assign addr[1324]= -76474970;
assign addr[1325]= -152852926;
assign addr[1326]= -229036977;
assign addr[1327]= -304930476;
assign addr[1328]= -380437148;
assign addr[1329]= -455461206;
assign addr[1330]= -529907477;
assign addr[1331]= -603681519;
assign addr[1332]= -676689746;
assign addr[1333]= -748839539;
assign addr[1334]= -820039373;
assign addr[1335]= -890198924;
assign addr[1336]= -959229189;
assign addr[1337]= -1027042599;
assign addr[1338]= -1093553126;
assign addr[1339]= -1158676398;
assign addr[1340]= -1222329801;
assign addr[1341]= -1284432584;
assign addr[1342]= -1344905966;
assign addr[1343]= -1403673233;
assign addr[1344]= -1460659832;
assign addr[1345]= -1515793473;
assign addr[1346]= -1569004214;
assign addr[1347]= -1620224553;
assign addr[1348]= -1669389513;
assign addr[1349]= -1716436725;
assign addr[1350]= -1761306505;
assign addr[1351]= -1803941934;
assign addr[1352]= -1844288924;
assign addr[1353]= -1882296293;
assign addr[1354]= -1917915825;
assign addr[1355]= -1951102334;
assign addr[1356]= -1981813720;
assign addr[1357]= -2010011024;
assign addr[1358]= -2035658475;
assign addr[1359]= -2058723538;
assign addr[1360]= -2079176953;
assign addr[1361]= -2096992772;
assign addr[1362]= -2112148396;
assign addr[1363]= -2124624598;
assign addr[1364]= -2134405552;
assign addr[1365]= -2141478848;
assign addr[1366]= -2145835515;
assign addr[1367]= -2147470025;
assign addr[1368]= -2146380306;
assign addr[1369]= -2142567738;
assign addr[1370]= -2136037160;
assign addr[1371]= -2126796855;
assign addr[1372]= -2114858546;
assign addr[1373]= -2100237377;
assign addr[1374]= -2082951896;
assign addr[1375]= -2063024031;
assign addr[1376]= -2040479063;
assign addr[1377]= -2015345591;
assign addr[1378]= -1987655498;
assign addr[1379]= -1957443913;
assign addr[1380]= -1924749160;
assign addr[1381]= -1889612716;
assign addr[1382]= -1852079154;
assign addr[1383]= -1812196087;
assign addr[1384]= -1770014111;
assign addr[1385]= -1725586737;
assign addr[1386]= -1678970324;
assign addr[1387]= -1630224009;
assign addr[1388]= -1579409630;
assign addr[1389]= -1526591649;
assign addr[1390]= -1471837070;
assign addr[1391]= -1415215352;
assign addr[1392]= -1356798326;
assign addr[1393]= -1296660098;
assign addr[1394]= -1234876957;
assign addr[1395]= -1171527280;
assign addr[1396]= -1106691431;
assign addr[1397]= -1040451659;
assign addr[1398]= -972891995;
assign addr[1399]= -904098143;
assign addr[1400]= -834157373;
assign addr[1401]= -763158411;
assign addr[1402]= -691191324;
assign addr[1403]= -618347408;
assign addr[1404]= -544719071;
assign addr[1405]= -470399716;
assign addr[1406]= -395483624;
assign addr[1407]= -320065829;
assign addr[1408]= -244242007;
assign addr[1409]= -168108346;
assign addr[1410]= -91761426;
assign addr[1411]= -15298099;
assign addr[1412]= 61184634;
assign addr[1413]= 137589750;
assign addr[1414]= 213820322;
assign addr[1415]= 289779648;
assign addr[1416]= 365371365;
assign addr[1417]= 440499581;
assign addr[1418]= 515068990;
assign addr[1419]= 588984994;
assign addr[1420]= 662153826;
assign addr[1421]= 734482665;
assign addr[1422]= 805879757;
assign addr[1423]= 876254528;
assign addr[1424]= 945517704;
assign addr[1425]= 1013581418;
assign addr[1426]= 1080359326;
assign addr[1427]= 1145766716;
assign addr[1428]= 1209720613;
assign addr[1429]= 1272139887;
assign addr[1430]= 1332945355;
assign addr[1431]= 1392059879;
assign addr[1432]= 1449408469;
assign addr[1433]= 1504918373;
assign addr[1434]= 1558519173;
assign addr[1435]= 1610142873;
assign addr[1436]= 1659723983;
assign addr[1437]= 1707199606;
assign addr[1438]= 1752509516;
assign addr[1439]= 1795596234;
assign addr[1440]= 1836405100;
assign addr[1441]= 1874884346;
assign addr[1442]= 1910985158;
assign addr[1443]= 1944661739;
assign addr[1444]= 1975871368;
assign addr[1445]= 2004574453;
assign addr[1446]= 2030734582;
assign addr[1447]= 2054318569;
assign addr[1448]= 2075296495;
assign addr[1449]= 2093641749;
assign addr[1450]= 2109331059;
assign addr[1451]= 2122344521;
assign addr[1452]= 2132665626;
assign addr[1453]= 2140281282;
assign addr[1454]= 2145181827;
assign addr[1455]= 2147361045;
assign addr[1456]= 2146816171;
assign addr[1457]= 2143547897;
assign addr[1458]= 2137560369;
assign addr[1459]= 2128861181;
assign addr[1460]= 2117461370;
assign addr[1461]= 2103375398;
assign addr[1462]= 2086621133;
assign addr[1463]= 2067219829;
assign addr[1464]= 2045196100;
assign addr[1465]= 2020577882;
assign addr[1466]= 1993396407;
assign addr[1467]= 1963686155;
assign addr[1468]= 1931484818;
assign addr[1469]= 1896833245;
assign addr[1470]= 1859775393;
assign addr[1471]= 1820358275;
assign addr[1472]= 1778631892;
assign addr[1473]= 1734649179;
assign addr[1474]= 1688465931;
assign addr[1475]= 1640140734;
assign addr[1476]= 1589734894;
assign addr[1477]= 1537312353;
assign addr[1478]= 1482939614;
assign addr[1479]= 1426685652;
assign addr[1480]= 1368621831;
assign addr[1481]= 1308821808;
assign addr[1482]= 1247361445;
assign addr[1483]= 1184318708;
assign addr[1484]= 1119773573;
assign addr[1485]= 1053807919;
assign addr[1486]= 986505429;
assign addr[1487]= 917951481;
assign addr[1488]= 848233042;
assign addr[1489]= 777438554;
assign addr[1490]= 705657826;
assign addr[1491]= 632981917;
assign addr[1492]= 559503022;
assign addr[1493]= 485314355;
assign addr[1494]= 410510029;
assign addr[1495]= 335184940;
assign addr[1496]= 259434643;
assign addr[1497]= 183355234;
assign addr[1498]= 107043224;
assign addr[1499]= 30595422;
assign addr[1500]= -45891193;
assign addr[1501]= -122319591;
assign addr[1502]= -198592817;
assign addr[1503]= -274614114;
assign addr[1504]= -350287041;
assign addr[1505]= -425515602;
assign addr[1506]= -500204365;
assign addr[1507]= -574258580;
assign addr[1508]= -647584304;
assign addr[1509]= -720088517;
assign addr[1510]= -791679244;
assign addr[1511]= -862265664;
assign addr[1512]= -931758235;
assign addr[1513]= -1000068799;
assign addr[1514]= -1067110699;
assign addr[1515]= -1132798888;
assign addr[1516]= -1197050035;
assign addr[1517]= -1259782632;
assign addr[1518]= -1320917099;
assign addr[1519]= -1380375881;
assign addr[1520]= -1438083551;
assign addr[1521]= -1493966902;
assign addr[1522]= -1547955041;
assign addr[1523]= -1599979481;
assign addr[1524]= -1649974225;
assign addr[1525]= -1697875851;
assign addr[1526]= -1743623590;
assign addr[1527]= -1787159411;
assign addr[1528]= -1828428082;
assign addr[1529]= -1867377253;
assign addr[1530]= -1903957513;
assign addr[1531]= -1938122457;
assign addr[1532]= -1969828744;
assign addr[1533]= -1999036154;
assign addr[1534]= -2025707632;
assign addr[1535]= -2049809346;
assign addr[1536]= -2071310720;
assign addr[1537]= -2090184478;
assign addr[1538]= -2106406677;
assign addr[1539]= -2119956737;
assign addr[1540]= -2130817471;
assign addr[1541]= -2138975100;
assign addr[1542]= -2144419275;
assign addr[1543]= -2147143090;
assign addr[1544]= -2147143090;
assign addr[1545]= -2144419275;
assign addr[1546]= -2138975100;
assign addr[1547]= -2130817471;
assign addr[1548]= -2119956737;
assign addr[1549]= -2106406677;
assign addr[1550]= -2090184478;
assign addr[1551]= -2071310720;
assign addr[1552]= -2049809346;
assign addr[1553]= -2025707632;
assign addr[1554]= -1999036154;
assign addr[1555]= -1969828744;
assign addr[1556]= -1938122457;
assign addr[1557]= -1903957513;
assign addr[1558]= -1867377253;
assign addr[1559]= -1828428082;
assign addr[1560]= -1787159411;
assign addr[1561]= -1743623590;
assign addr[1562]= -1697875851;
assign addr[1563]= -1649974225;
assign addr[1564]= -1599979481;
assign addr[1565]= -1547955041;
assign addr[1566]= -1493966902;
assign addr[1567]= -1438083551;
assign addr[1568]= -1380375881;
assign addr[1569]= -1320917099;
assign addr[1570]= -1259782632;
assign addr[1571]= -1197050035;
assign addr[1572]= -1132798888;
assign addr[1573]= -1067110699;
assign addr[1574]= -1000068799;
assign addr[1575]= -931758235;
assign addr[1576]= -862265664;
assign addr[1577]= -791679244;
assign addr[1578]= -720088517;
assign addr[1579]= -647584304;
assign addr[1580]= -574258580;
assign addr[1581]= -500204365;
assign addr[1582]= -425515602;
assign addr[1583]= -350287041;
assign addr[1584]= -274614114;
assign addr[1585]= -198592817;
assign addr[1586]= -122319591;
assign addr[1587]= -45891193;
assign addr[1588]= 30595422;
assign addr[1589]= 107043224;
assign addr[1590]= 183355234;
assign addr[1591]= 259434643;
assign addr[1592]= 335184940;
assign addr[1593]= 410510029;
assign addr[1594]= 485314355;
assign addr[1595]= 559503022;
assign addr[1596]= 632981917;
assign addr[1597]= 705657826;
assign addr[1598]= 777438554;
assign addr[1599]= 848233042;
assign addr[1600]= 917951481;
assign addr[1601]= 986505429;
assign addr[1602]= 1053807919;
assign addr[1603]= 1119773573;
assign addr[1604]= 1184318708;
assign addr[1605]= 1247361445;
assign addr[1606]= 1308821808;
assign addr[1607]= 1368621831;
assign addr[1608]= 1426685652;
assign addr[1609]= 1482939614;
assign addr[1610]= 1537312353;
assign addr[1611]= 1589734894;
assign addr[1612]= 1640140734;
assign addr[1613]= 1688465931;
assign addr[1614]= 1734649179;
assign addr[1615]= 1778631892;
assign addr[1616]= 1820358275;
assign addr[1617]= 1859775393;
assign addr[1618]= 1896833245;
assign addr[1619]= 1931484818;
assign addr[1620]= 1963686155;
assign addr[1621]= 1993396407;
assign addr[1622]= 2020577882;
assign addr[1623]= 2045196100;
assign addr[1624]= 2067219829;
assign addr[1625]= 2086621133;
assign addr[1626]= 2103375398;
assign addr[1627]= 2117461370;
assign addr[1628]= 2128861181;
assign addr[1629]= 2137560369;
assign addr[1630]= 2143547897;
assign addr[1631]= 2146816171;
assign addr[1632]= 2147361045;
assign addr[1633]= 2145181827;
assign addr[1634]= 2140281282;
assign addr[1635]= 2132665626;
assign addr[1636]= 2122344521;
assign addr[1637]= 2109331059;
assign addr[1638]= 2093641749;
assign addr[1639]= 2075296495;
assign addr[1640]= 2054318569;
assign addr[1641]= 2030734582;
assign addr[1642]= 2004574453;
assign addr[1643]= 1975871368;
assign addr[1644]= 1944661739;
assign addr[1645]= 1910985158;
assign addr[1646]= 1874884346;
assign addr[1647]= 1836405100;
assign addr[1648]= 1795596234;
assign addr[1649]= 1752509516;
assign addr[1650]= 1707199606;
assign addr[1651]= 1659723983;
assign addr[1652]= 1610142873;
assign addr[1653]= 1558519173;
assign addr[1654]= 1504918373;
assign addr[1655]= 1449408469;
assign addr[1656]= 1392059879;
assign addr[1657]= 1332945355;
assign addr[1658]= 1272139887;
assign addr[1659]= 1209720613;
assign addr[1660]= 1145766716;
assign addr[1661]= 1080359326;
assign addr[1662]= 1013581418;
assign addr[1663]= 945517704;
assign addr[1664]= 876254528;
assign addr[1665]= 805879757;
assign addr[1666]= 734482665;
assign addr[1667]= 662153826;
assign addr[1668]= 588984994;
assign addr[1669]= 515068990;
assign addr[1670]= 440499581;
assign addr[1671]= 365371365;
assign addr[1672]= 289779648;
assign addr[1673]= 213820322;
assign addr[1674]= 137589750;
assign addr[1675]= 61184634;
assign addr[1676]= -15298099;
assign addr[1677]= -91761426;
assign addr[1678]= -168108346;
assign addr[1679]= -244242007;
assign addr[1680]= -320065829;
assign addr[1681]= -395483624;
assign addr[1682]= -470399716;
assign addr[1683]= -544719071;
assign addr[1684]= -618347408;
assign addr[1685]= -691191324;
assign addr[1686]= -763158411;
assign addr[1687]= -834157373;
assign addr[1688]= -904098143;
assign addr[1689]= -972891995;
assign addr[1690]= -1040451659;
assign addr[1691]= -1106691431;
assign addr[1692]= -1171527280;
assign addr[1693]= -1234876957;
assign addr[1694]= -1296660098;
assign addr[1695]= -1356798326;
assign addr[1696]= -1415215352;
assign addr[1697]= -1471837070;
assign addr[1698]= -1526591649;
assign addr[1699]= -1579409630;
assign addr[1700]= -1630224009;
assign addr[1701]= -1678970324;
assign addr[1702]= -1725586737;
assign addr[1703]= -1770014111;
assign addr[1704]= -1812196087;
assign addr[1705]= -1852079154;
assign addr[1706]= -1889612716;
assign addr[1707]= -1924749160;
assign addr[1708]= -1957443913;
assign addr[1709]= -1987655498;
assign addr[1710]= -2015345591;
assign addr[1711]= -2040479063;
assign addr[1712]= -2063024031;
assign addr[1713]= -2082951896;
assign addr[1714]= -2100237377;
assign addr[1715]= -2114858546;
assign addr[1716]= -2126796855;
assign addr[1717]= -2136037160;
assign addr[1718]= -2142567738;
assign addr[1719]= -2146380306;
assign addr[1720]= -2147470025;
assign addr[1721]= -2145835515;
assign addr[1722]= -2141478848;
assign addr[1723]= -2134405552;
assign addr[1724]= -2124624598;
assign addr[1725]= -2112148396;
assign addr[1726]= -2096992772;
assign addr[1727]= -2079176953;
assign addr[1728]= -2058723538;
assign addr[1729]= -2035658475;
assign addr[1730]= -2010011024;
assign addr[1731]= -1981813720;
assign addr[1732]= -1951102334;
assign addr[1733]= -1917915825;
assign addr[1734]= -1882296293;
assign addr[1735]= -1844288924;
assign addr[1736]= -1803941934;
assign addr[1737]= -1761306505;
assign addr[1738]= -1716436725;
assign addr[1739]= -1669389513;
assign addr[1740]= -1620224553;
assign addr[1741]= -1569004214;
assign addr[1742]= -1515793473;
assign addr[1743]= -1460659832;
assign addr[1744]= -1403673233;
assign addr[1745]= -1344905966;
assign addr[1746]= -1284432584;
assign addr[1747]= -1222329801;
assign addr[1748]= -1158676398;
assign addr[1749]= -1093553126;
assign addr[1750]= -1027042599;
assign addr[1751]= -959229189;
assign addr[1752]= -890198924;
assign addr[1753]= -820039373;
assign addr[1754]= -748839539;
assign addr[1755]= -676689746;
assign addr[1756]= -603681519;
assign addr[1757]= -529907477;
assign addr[1758]= -455461206;
assign addr[1759]= -380437148;
assign addr[1760]= -304930476;
assign addr[1761]= -229036977;
assign addr[1762]= -152852926;
assign addr[1763]= -76474970;
assign addr[1764]= 0;
assign addr[1765]= 76474970;
assign addr[1766]= 152852926;
assign addr[1767]= 229036977;
assign addr[1768]= 304930476;
assign addr[1769]= 380437148;
assign addr[1770]= 455461206;
assign addr[1771]= 529907477;
assign addr[1772]= 603681519;
assign addr[1773]= 676689746;
assign addr[1774]= 748839539;
assign addr[1775]= 820039373;
assign addr[1776]= 890198924;
assign addr[1777]= 959229189;
assign addr[1778]= 1027042599;
assign addr[1779]= 1093553126;
assign addr[1780]= 1158676398;
assign addr[1781]= 1222329801;
assign addr[1782]= 1284432584;
assign addr[1783]= 1344905966;
assign addr[1784]= 1403673233;
assign addr[1785]= 1460659832;
assign addr[1786]= 1515793473;
assign addr[1787]= 1569004214;
assign addr[1788]= 1620224553;
assign addr[1789]= 1669389513;
assign addr[1790]= 1716436725;
assign addr[1791]= 1761306505;
assign addr[1792]= 1803941934;
assign addr[1793]= 1844288924;
assign addr[1794]= 1882296293;
assign addr[1795]= 1917915825;
assign addr[1796]= 1951102334;
assign addr[1797]= 1981813720;
assign addr[1798]= 2010011024;
assign addr[1799]= 2035658475;
assign addr[1800]= 2058723538;
assign addr[1801]= 2079176953;
assign addr[1802]= 2096992772;
assign addr[1803]= 2112148396;
assign addr[1804]= 2124624598;
assign addr[1805]= 2134405552;
assign addr[1806]= 2141478848;
assign addr[1807]= 2145835515;
assign addr[1808]= 2147470025;
assign addr[1809]= 2146380306;
assign addr[1810]= 2142567738;
assign addr[1811]= 2136037160;
assign addr[1812]= 2126796855;
assign addr[1813]= 2114858546;
assign addr[1814]= 2100237377;
assign addr[1815]= 2082951896;
assign addr[1816]= 2063024031;
assign addr[1817]= 2040479063;
assign addr[1818]= 2015345591;
assign addr[1819]= 1987655498;
assign addr[1820]= 1957443913;
assign addr[1821]= 1924749160;
assign addr[1822]= 1889612716;
assign addr[1823]= 1852079154;
assign addr[1824]= 1812196087;
assign addr[1825]= 1770014111;
assign addr[1826]= 1725586737;
assign addr[1827]= 1678970324;
assign addr[1828]= 1630224009;
assign addr[1829]= 1579409630;
assign addr[1830]= 1526591649;
assign addr[1831]= 1471837070;
assign addr[1832]= 1415215352;
assign addr[1833]= 1356798326;
assign addr[1834]= 1296660098;
assign addr[1835]= 1234876957;
assign addr[1836]= 1171527280;
assign addr[1837]= 1106691431;
assign addr[1838]= 1040451659;
assign addr[1839]= 972891995;
assign addr[1840]= 904098143;
assign addr[1841]= 834157373;
assign addr[1842]= 763158411;
assign addr[1843]= 691191324;
assign addr[1844]= 618347408;
assign addr[1845]= 544719071;
assign addr[1846]= 470399716;
assign addr[1847]= 395483624;
assign addr[1848]= 320065829;
assign addr[1849]= 244242007;
assign addr[1850]= 168108346;
assign addr[1851]= 91761426;
assign addr[1852]= 15298099;
assign addr[1853]= -61184634;
assign addr[1854]= -137589750;
assign addr[1855]= -213820322;
assign addr[1856]= -289779648;
assign addr[1857]= -365371365;
assign addr[1858]= -440499581;
assign addr[1859]= -515068990;
assign addr[1860]= -588984994;
assign addr[1861]= -662153826;
assign addr[1862]= -734482665;
assign addr[1863]= -805879757;
assign addr[1864]= -876254528;
assign addr[1865]= -945517704;
assign addr[1866]= -1013581418;
assign addr[1867]= -1080359326;
assign addr[1868]= -1145766716;
assign addr[1869]= -1209720613;
assign addr[1870]= -1272139887;
assign addr[1871]= -1332945355;
assign addr[1872]= -1392059879;
assign addr[1873]= -1449408469;
assign addr[1874]= -1504918373;
assign addr[1875]= -1558519173;
assign addr[1876]= -1610142873;
assign addr[1877]= -1659723983;
assign addr[1878]= -1707199606;
assign addr[1879]= -1752509516;
assign addr[1880]= -1795596234;
assign addr[1881]= -1836405100;
assign addr[1882]= -1874884346;
assign addr[1883]= -1910985158;
assign addr[1884]= -1944661739;
assign addr[1885]= -1975871368;
assign addr[1886]= -2004574453;
assign addr[1887]= -2030734582;
assign addr[1888]= -2054318569;
assign addr[1889]= -2075296495;
assign addr[1890]= -2093641749;
assign addr[1891]= -2109331059;
assign addr[1892]= -2122344521;
assign addr[1893]= -2132665626;
assign addr[1894]= -2140281282;
assign addr[1895]= -2145181827;
assign addr[1896]= -2147361045;
assign addr[1897]= -2146816171;
assign addr[1898]= -2143547897;
assign addr[1899]= -2137560369;
assign addr[1900]= -2128861181;
assign addr[1901]= -2117461370;
assign addr[1902]= -2103375398;
assign addr[1903]= -2086621133;
assign addr[1904]= -2067219829;
assign addr[1905]= -2045196100;
assign addr[1906]= -2020577882;
assign addr[1907]= -1993396407;
assign addr[1908]= -1963686155;
assign addr[1909]= -1931484818;
assign addr[1910]= -1896833245;
assign addr[1911]= -1859775393;
assign addr[1912]= -1820358275;
assign addr[1913]= -1778631892;
assign addr[1914]= -1734649179;
assign addr[1915]= -1688465931;
assign addr[1916]= -1640140734;
assign addr[1917]= -1589734894;
assign addr[1918]= -1537312353;
assign addr[1919]= -1482939614;
assign addr[1920]= -1426685652;
assign addr[1921]= -1368621831;
assign addr[1922]= -1308821808;
assign addr[1923]= -1247361445;
assign addr[1924]= -1184318708;
assign addr[1925]= -1119773573;
assign addr[1926]= -1053807919;
assign addr[1927]= -986505429;
assign addr[1928]= -917951481;
assign addr[1929]= -848233042;
assign addr[1930]= -777438554;
assign addr[1931]= -705657826;
assign addr[1932]= -632981917;
assign addr[1933]= -559503022;
assign addr[1934]= -485314355;
assign addr[1935]= -410510029;
assign addr[1936]= -335184940;
assign addr[1937]= -259434643;
assign addr[1938]= -183355234;
assign addr[1939]= -107043224;
assign addr[1940]= -30595422;
assign addr[1941]= 45891193;
assign addr[1942]= 122319591;
assign addr[1943]= 198592817;
assign addr[1944]= 274614114;
assign addr[1945]= 350287041;
assign addr[1946]= 425515602;
assign addr[1947]= 500204365;
assign addr[1948]= 574258580;
assign addr[1949]= 647584304;
assign addr[1950]= 720088517;
assign addr[1951]= 791679244;
assign addr[1952]= 862265664;
assign addr[1953]= 931758235;
assign addr[1954]= 1000068799;
assign addr[1955]= 1067110699;
assign addr[1956]= 1132798888;
assign addr[1957]= 1197050035;
assign addr[1958]= 1259782632;
assign addr[1959]= 1320917099;
assign addr[1960]= 1380375881;
assign addr[1961]= 1438083551;
assign addr[1962]= 1493966902;
assign addr[1963]= 1547955041;
assign addr[1964]= 1599979481;
assign addr[1965]= 1649974225;
assign addr[1966]= 1697875851;
assign addr[1967]= 1743623590;
assign addr[1968]= 1787159411;
assign addr[1969]= 1828428082;
assign addr[1970]= 1867377253;
assign addr[1971]= 1903957513;
assign addr[1972]= 1938122457;
assign addr[1973]= 1969828744;
assign addr[1974]= 1999036154;
assign addr[1975]= 2025707632;
assign addr[1976]= 2049809346;
assign addr[1977]= 2071310720;
assign addr[1978]= 2090184478;
assign addr[1979]= 2106406677;
assign addr[1980]= 2119956737;
assign addr[1981]= 2130817471;
assign addr[1982]= 2138975100;
assign addr[1983]= 2144419275;
assign addr[1984]= 2147143090;
assign addr[1985]= 2147143090;
assign addr[1986]= 2144419275;
assign addr[1987]= 2138975100;
assign addr[1988]= 2130817471;
assign addr[1989]= 2119956737;
assign addr[1990]= 2106406677;
assign addr[1991]= 2090184478;
assign addr[1992]= 2071310720;
assign addr[1993]= 2049809346;
assign addr[1994]= 2025707632;
assign addr[1995]= 1999036154;
assign addr[1996]= 1969828744;
assign addr[1997]= 1938122457;
assign addr[1998]= 1903957513;
assign addr[1999]= 1867377253;
assign addr[2000]= 1828428082;
assign addr[2001]= 1787159411;
assign addr[2002]= 1743623590;
assign addr[2003]= 1697875851;
assign addr[2004]= 1649974225;
assign addr[2005]= 1599979481;
assign addr[2006]= 1547955041;
assign addr[2007]= 1493966902;
assign addr[2008]= 1438083551;
assign addr[2009]= 1380375881;
assign addr[2010]= 1320917099;
assign addr[2011]= 1259782632;
assign addr[2012]= 1197050035;
assign addr[2013]= 1132798888;
assign addr[2014]= 1067110699;
assign addr[2015]= 1000068799;
assign addr[2016]= 931758235;
assign addr[2017]= 862265664;
assign addr[2018]= 791679244;
assign addr[2019]= 720088517;
assign addr[2020]= 647584304;
assign addr[2021]= 574258580;
assign addr[2022]= 500204365;
assign addr[2023]= 425515602;
assign addr[2024]= 350287041;
assign addr[2025]= 274614114;
assign addr[2026]= 198592817;
assign addr[2027]= 122319591;
assign addr[2028]= 45891193;
assign addr[2029]= -30595422;
assign addr[2030]= -107043224;
assign addr[2031]= -183355234;
assign addr[2032]= -259434643;
assign addr[2033]= -335184940;
assign addr[2034]= -410510029;
assign addr[2035]= -485314355;
assign addr[2036]= -559503022;
assign addr[2037]= -632981917;
assign addr[2038]= -705657826;
assign addr[2039]= -777438554;
assign addr[2040]= -848233042;
assign addr[2041]= -917951481;
assign addr[2042]= -986505429;
assign addr[2043]= -1053807919;
assign addr[2044]= -1119773573;
assign addr[2045]= -1184318708;
assign addr[2046]= -1247361445;
assign addr[2047]= -1308821808;
assign addr[2048]= -1368621831;
assign addr[2049]= -1426685652;
assign addr[2050]= -1482939614;
assign addr[2051]= -1537312353;
assign addr[2052]= -1589734894;
assign addr[2053]= -1640140734;
assign addr[2054]= -1688465931;
assign addr[2055]= -1734649179;
assign addr[2056]= -1778631892;
assign addr[2057]= -1820358275;
assign addr[2058]= -1859775393;
assign addr[2059]= -1896833245;
assign addr[2060]= -1931484818;
assign addr[2061]= -1963686155;
assign addr[2062]= -1993396407;
assign addr[2063]= -2020577882;
assign addr[2064]= -2045196100;
assign addr[2065]= -2067219829;
assign addr[2066]= -2086621133;
assign addr[2067]= -2103375398;
assign addr[2068]= -2117461370;
assign addr[2069]= -2128861181;
assign addr[2070]= -2137560369;
assign addr[2071]= -2143547897;
assign addr[2072]= -2146816171;
assign addr[2073]= -2147361045;
assign addr[2074]= -2145181827;
assign addr[2075]= -2140281282;
assign addr[2076]= -2132665626;
assign addr[2077]= -2122344521;
assign addr[2078]= -2109331059;
assign addr[2079]= -2093641749;
assign addr[2080]= -2075296495;
assign addr[2081]= -2054318569;
assign addr[2082]= -2030734582;
assign addr[2083]= -2004574453;
assign addr[2084]= -1975871368;
assign addr[2085]= -1944661739;
assign addr[2086]= -1910985158;
assign addr[2087]= -1874884346;
assign addr[2088]= -1836405100;
assign addr[2089]= -1795596234;
assign addr[2090]= -1752509516;
assign addr[2091]= -1707199606;
assign addr[2092]= -1659723983;
assign addr[2093]= -1610142873;
assign addr[2094]= -1558519173;
assign addr[2095]= -1504918373;
assign addr[2096]= -1449408469;
assign addr[2097]= -1392059879;
assign addr[2098]= -1332945355;
assign addr[2099]= -1272139887;
assign addr[2100]= -1209720613;
assign addr[2101]= -1145766716;
assign addr[2102]= -1080359326;
assign addr[2103]= -1013581418;
assign addr[2104]= -945517704;
assign addr[2105]= -876254528;
assign addr[2106]= -805879757;
assign addr[2107]= -734482665;
assign addr[2108]= -662153826;
assign addr[2109]= -588984994;
assign addr[2110]= -515068990;
assign addr[2111]= -440499581;
assign addr[2112]= -365371365;
assign addr[2113]= -289779648;
assign addr[2114]= -213820322;
assign addr[2115]= -137589750;
assign addr[2116]= -61184634;
assign addr[2117]= 15298099;
assign addr[2118]= 91761426;
assign addr[2119]= 168108346;
assign addr[2120]= 244242007;
assign addr[2121]= 320065829;
assign addr[2122]= 395483624;
assign addr[2123]= 470399716;
assign addr[2124]= 544719071;
assign addr[2125]= 618347408;
assign addr[2126]= 691191324;
assign addr[2127]= 763158411;
assign addr[2128]= 834157373;
assign addr[2129]= 904098143;
assign addr[2130]= 972891995;
assign addr[2131]= 1040451659;
assign addr[2132]= 1106691431;
assign addr[2133]= 1171527280;
assign addr[2134]= 1234876957;
assign addr[2135]= 1296660098;
assign addr[2136]= 1356798326;
assign addr[2137]= 1415215352;
assign addr[2138]= 1471837070;
assign addr[2139]= 1526591649;
assign addr[2140]= 1579409630;
assign addr[2141]= 1630224009;
assign addr[2142]= 1678970324;
assign addr[2143]= 1725586737;
assign addr[2144]= 1770014111;
assign addr[2145]= 1812196087;
assign addr[2146]= 1852079154;
assign addr[2147]= 1889612716;
assign addr[2148]= 1924749160;
assign addr[2149]= 1957443913;
assign addr[2150]= 1987655498;
assign addr[2151]= 2015345591;
assign addr[2152]= 2040479063;
assign addr[2153]= 2063024031;
assign addr[2154]= 2082951896;
assign addr[2155]= 2100237377;
assign addr[2156]= 2114858546;
assign addr[2157]= 2126796855;
assign addr[2158]= 2136037160;
assign addr[2159]= 2142567738;
assign addr[2160]= 2146380306;
assign addr[2161]= 2147470025;
assign addr[2162]= 2145835515;
assign addr[2163]= 2141478848;
assign addr[2164]= 2134405552;
assign addr[2165]= 2124624598;
assign addr[2166]= 2112148396;
assign addr[2167]= 2096992772;
assign addr[2168]= 2079176953;
assign addr[2169]= 2058723538;
assign addr[2170]= 2035658475;
assign addr[2171]= 2010011024;
assign addr[2172]= 1981813720;
assign addr[2173]= 1951102334;
assign addr[2174]= 1917915825;
assign addr[2175]= 1882296293;
assign addr[2176]= 1844288924;
assign addr[2177]= 1803941934;
assign addr[2178]= 1761306505;
assign addr[2179]= 1716436725;
assign addr[2180]= 1669389513;
assign addr[2181]= 1620224553;
assign addr[2182]= 1569004214;
assign addr[2183]= 1515793473;
assign addr[2184]= 1460659832;
assign addr[2185]= 1403673233;
assign addr[2186]= 1344905966;
assign addr[2187]= 1284432584;
assign addr[2188]= 1222329801;
assign addr[2189]= 1158676398;
assign addr[2190]= 1093553126;
assign addr[2191]= 1027042599;
assign addr[2192]= 959229189;
assign addr[2193]= 890198924;
assign addr[2194]= 820039373;
assign addr[2195]= 748839539;
assign addr[2196]= 676689746;
assign addr[2197]= 603681519;
assign addr[2198]= 529907477;
assign addr[2199]= 455461206;
assign addr[2200]= 380437148;
assign addr[2201]= 304930476;
assign addr[2202]= 229036977;
assign addr[2203]= 152852926;
assign addr[2204]= 76474970;
assign addr[2205]= 0;
assign addr[2206]= -76474970;
assign addr[2207]= -152852926;
assign addr[2208]= -229036977;
assign addr[2209]= -304930476;
assign addr[2210]= -380437148;
assign addr[2211]= -455461206;
assign addr[2212]= -529907477;
assign addr[2213]= -603681519;
assign addr[2214]= -676689746;
assign addr[2215]= -748839539;
assign addr[2216]= -820039373;
assign addr[2217]= -890198924;
assign addr[2218]= -959229189;
assign addr[2219]= -1027042599;
assign addr[2220]= -1093553126;
assign addr[2221]= -1158676398;
assign addr[2222]= -1222329801;
assign addr[2223]= -1284432584;
assign addr[2224]= -1344905966;
assign addr[2225]= -1403673233;
assign addr[2226]= -1460659832;
assign addr[2227]= -1515793473;
assign addr[2228]= -1569004214;
assign addr[2229]= -1620224553;
assign addr[2230]= -1669389513;
assign addr[2231]= -1716436725;
assign addr[2232]= -1761306505;
assign addr[2233]= -1803941934;
assign addr[2234]= -1844288924;
assign addr[2235]= -1882296293;
assign addr[2236]= -1917915825;
assign addr[2237]= -1951102334;
assign addr[2238]= -1981813720;
assign addr[2239]= -2010011024;
assign addr[2240]= -2035658475;
assign addr[2241]= -2058723538;
assign addr[2242]= -2079176953;
assign addr[2243]= -2096992772;
assign addr[2244]= -2112148396;
assign addr[2245]= -2124624598;
assign addr[2246]= -2134405552;
assign addr[2247]= -2141478848;
assign addr[2248]= -2145835515;
assign addr[2249]= -2147470025;
assign addr[2250]= -2146380306;
assign addr[2251]= -2142567738;
assign addr[2252]= -2136037160;
assign addr[2253]= -2126796855;
assign addr[2254]= -2114858546;
assign addr[2255]= -2100237377;
assign addr[2256]= -2082951896;
assign addr[2257]= -2063024031;
assign addr[2258]= -2040479063;
assign addr[2259]= -2015345591;
assign addr[2260]= -1987655498;
assign addr[2261]= -1957443913;
assign addr[2262]= -1924749160;
assign addr[2263]= -1889612716;
assign addr[2264]= -1852079154;
assign addr[2265]= -1812196087;
assign addr[2266]= -1770014111;
assign addr[2267]= -1725586737;
assign addr[2268]= -1678970324;
assign addr[2269]= -1630224009;
assign addr[2270]= -1579409630;
assign addr[2271]= -1526591649;
assign addr[2272]= -1471837070;
assign addr[2273]= -1415215352;
assign addr[2274]= -1356798326;
assign addr[2275]= -1296660098;
assign addr[2276]= -1234876957;
assign addr[2277]= -1171527280;
assign addr[2278]= -1106691431;
assign addr[2279]= -1040451659;
assign addr[2280]= -972891995;
assign addr[2281]= -904098143;
assign addr[2282]= -834157373;
assign addr[2283]= -763158411;
assign addr[2284]= -691191324;
assign addr[2285]= -618347408;
assign addr[2286]= -544719071;
assign addr[2287]= -470399716;
assign addr[2288]= -395483624;
assign addr[2289]= -320065829;
assign addr[2290]= -244242007;
assign addr[2291]= -168108346;
assign addr[2292]= -91761426;
assign addr[2293]= -15298099;
assign addr[2294]= 61184634;
assign addr[2295]= 137589750;
assign addr[2296]= 213820322;
assign addr[2297]= 289779648;
assign addr[2298]= 365371365;
assign addr[2299]= 440499581;
assign addr[2300]= 515068990;
assign addr[2301]= 588984994;
assign addr[2302]= 662153826;
assign addr[2303]= 734482665;
assign addr[2304]= 805879757;
assign addr[2305]= 876254528;
assign addr[2306]= 945517704;
assign addr[2307]= 1013581418;
assign addr[2308]= 1080359326;
assign addr[2309]= 1145766716;
assign addr[2310]= 1209720613;
assign addr[2311]= 1272139887;
assign addr[2312]= 1332945355;
assign addr[2313]= 1392059879;
assign addr[2314]= 1449408469;
assign addr[2315]= 1504918373;
assign addr[2316]= 1558519173;
assign addr[2317]= 1610142873;
assign addr[2318]= 1659723983;
assign addr[2319]= 1707199606;
assign addr[2320]= 1752509516;
assign addr[2321]= 1795596234;
assign addr[2322]= 1836405100;
assign addr[2323]= 1874884346;
assign addr[2324]= 1910985158;
assign addr[2325]= 1944661739;
assign addr[2326]= 1975871368;
assign addr[2327]= 2004574453;
assign addr[2328]= 2030734582;
assign addr[2329]= 2054318569;
assign addr[2330]= 2075296495;
assign addr[2331]= 2093641749;
assign addr[2332]= 2109331059;
assign addr[2333]= 2122344521;
assign addr[2334]= 2132665626;
assign addr[2335]= 2140281282;
assign addr[2336]= 2145181827;
assign addr[2337]= 2147361045;
assign addr[2338]= 2146816171;
assign addr[2339]= 2143547897;
assign addr[2340]= 2137560369;
assign addr[2341]= 2128861181;
assign addr[2342]= 2117461370;
assign addr[2343]= 2103375398;
assign addr[2344]= 2086621133;
assign addr[2345]= 2067219829;
assign addr[2346]= 2045196100;
assign addr[2347]= 2020577882;
assign addr[2348]= 1993396407;
assign addr[2349]= 1963686155;
assign addr[2350]= 1931484818;
assign addr[2351]= 1896833245;
assign addr[2352]= 1859775393;
assign addr[2353]= 1820358275;
assign addr[2354]= 1778631892;
assign addr[2355]= 1734649179;
assign addr[2356]= 1688465931;
assign addr[2357]= 1640140734;
assign addr[2358]= 1589734894;
assign addr[2359]= 1537312353;
assign addr[2360]= 1482939614;
assign addr[2361]= 1426685652;
assign addr[2362]= 1368621831;
assign addr[2363]= 1308821808;
assign addr[2364]= 1247361445;
assign addr[2365]= 1184318708;
assign addr[2366]= 1119773573;
assign addr[2367]= 1053807919;
assign addr[2368]= 986505429;
assign addr[2369]= 917951481;
assign addr[2370]= 848233042;
assign addr[2371]= 777438554;
assign addr[2372]= 705657826;
assign addr[2373]= 632981917;
assign addr[2374]= 559503022;
assign addr[2375]= 485314355;
assign addr[2376]= 410510029;
assign addr[2377]= 335184940;
assign addr[2378]= 259434643;
assign addr[2379]= 183355234;
assign addr[2380]= 107043224;
assign addr[2381]= 30595422;
assign addr[2382]= -45891193;
assign addr[2383]= -122319591;
assign addr[2384]= -198592817;
assign addr[2385]= -274614114;
assign addr[2386]= -350287041;
assign addr[2387]= -425515602;
assign addr[2388]= -500204365;
assign addr[2389]= -574258580;
assign addr[2390]= -647584304;
assign addr[2391]= -720088517;
assign addr[2392]= -791679244;
assign addr[2393]= -862265664;
assign addr[2394]= -931758235;
assign addr[2395]= -1000068799;
assign addr[2396]= -1067110699;
assign addr[2397]= -1132798888;
assign addr[2398]= -1197050035;
assign addr[2399]= -1259782632;
assign addr[2400]= -1320917099;
assign addr[2401]= -1380375881;
assign addr[2402]= -1438083551;
assign addr[2403]= -1493966902;
assign addr[2404]= -1547955041;
assign addr[2405]= -1599979481;
assign addr[2406]= -1649974225;
assign addr[2407]= -1697875851;
assign addr[2408]= -1743623590;
assign addr[2409]= -1787159411;
assign addr[2410]= -1828428082;
assign addr[2411]= -1867377253;
assign addr[2412]= -1903957513;
assign addr[2413]= -1938122457;
assign addr[2414]= -1969828744;
assign addr[2415]= -1999036154;
assign addr[2416]= -2025707632;
assign addr[2417]= -2049809346;
assign addr[2418]= -2071310720;
assign addr[2419]= -2090184478;
assign addr[2420]= -2106406677;
assign addr[2421]= -2119956737;
assign addr[2422]= -2130817471;
assign addr[2423]= -2138975100;
assign addr[2424]= -2144419275;
assign addr[2425]= -2147143090;
assign addr[2426]= -2147143090;
assign addr[2427]= -2144419275;
assign addr[2428]= -2138975100;
assign addr[2429]= -2130817471;
assign addr[2430]= -2119956737;
assign addr[2431]= -2106406677;
assign addr[2432]= -2090184478;
assign addr[2433]= -2071310720;
assign addr[2434]= -2049809346;
assign addr[2435]= -2025707632;
assign addr[2436]= -1999036154;
assign addr[2437]= -1969828744;
assign addr[2438]= -1938122457;
assign addr[2439]= -1903957513;
assign addr[2440]= -1867377253;
assign addr[2441]= -1828428082;
assign addr[2442]= -1787159411;
assign addr[2443]= -1743623590;
assign addr[2444]= -1697875851;
assign addr[2445]= -1649974225;
assign addr[2446]= -1599979481;
assign addr[2447]= -1547955041;
assign addr[2448]= -1493966902;
assign addr[2449]= -1438083551;
assign addr[2450]= -1380375881;
assign addr[2451]= -1320917099;
assign addr[2452]= -1259782632;
assign addr[2453]= -1197050035;
assign addr[2454]= -1132798888;
assign addr[2455]= -1067110699;
assign addr[2456]= -1000068799;
assign addr[2457]= -931758235;
assign addr[2458]= -862265664;
assign addr[2459]= -791679244;
assign addr[2460]= -720088517;
assign addr[2461]= -647584304;
assign addr[2462]= -574258580;
assign addr[2463]= -500204365;
assign addr[2464]= -425515602;
assign addr[2465]= -350287041;
assign addr[2466]= -274614114;
assign addr[2467]= -198592817;
assign addr[2468]= -122319591;
assign addr[2469]= -45891193;
assign addr[2470]= 30595422;
assign addr[2471]= 107043224;
assign addr[2472]= 183355234;
assign addr[2473]= 259434643;
assign addr[2474]= 335184940;
assign addr[2475]= 410510029;
assign addr[2476]= 485314355;
assign addr[2477]= 559503022;
assign addr[2478]= 632981917;
assign addr[2479]= 705657826;
assign addr[2480]= 777438554;
assign addr[2481]= 848233042;
assign addr[2482]= 917951481;
assign addr[2483]= 986505429;
assign addr[2484]= 1053807919;
assign addr[2485]= 1119773573;
assign addr[2486]= 1184318708;
assign addr[2487]= 1247361445;
assign addr[2488]= 1308821808;
assign addr[2489]= 1368621831;
assign addr[2490]= 1426685652;
assign addr[2491]= 1482939614;
assign addr[2492]= 1537312353;
assign addr[2493]= 1589734894;
assign addr[2494]= 1640140734;
assign addr[2495]= 1688465931;
assign addr[2496]= 1734649179;
assign addr[2497]= 1778631892;
assign addr[2498]= 1820358275;
assign addr[2499]= 1859775393;
assign addr[2500]= 1896833245;
assign addr[2501]= 1931484818;
assign addr[2502]= 1963686155;
assign addr[2503]= 1993396407;
assign addr[2504]= 2020577882;
assign addr[2505]= 2045196100;
assign addr[2506]= 2067219829;
assign addr[2507]= 2086621133;
assign addr[2508]= 2103375398;
assign addr[2509]= 2117461370;
assign addr[2510]= 2128861181;
assign addr[2511]= 2137560369;
assign addr[2512]= 2143547897;
assign addr[2513]= 2146816171;
assign addr[2514]= 2147361045;
assign addr[2515]= 2145181827;
assign addr[2516]= 2140281282;
assign addr[2517]= 2132665626;
assign addr[2518]= 2122344521;
assign addr[2519]= 2109331059;
assign addr[2520]= 2093641749;
assign addr[2521]= 2075296495;
assign addr[2522]= 2054318569;
assign addr[2523]= 2030734582;
assign addr[2524]= 2004574453;
assign addr[2525]= 1975871368;
assign addr[2526]= 1944661739;
assign addr[2527]= 1910985158;
assign addr[2528]= 1874884346;
assign addr[2529]= 1836405100;
assign addr[2530]= 1795596234;
assign addr[2531]= 1752509516;
assign addr[2532]= 1707199606;
assign addr[2533]= 1659723983;
assign addr[2534]= 1610142873;
assign addr[2535]= 1558519173;
assign addr[2536]= 1504918373;
assign addr[2537]= 1449408469;
assign addr[2538]= 1392059879;
assign addr[2539]= 1332945355;
assign addr[2540]= 1272139887;
assign addr[2541]= 1209720613;
assign addr[2542]= 1145766716;
assign addr[2543]= 1080359326;
assign addr[2544]= 1013581418;
assign addr[2545]= 945517704;
assign addr[2546]= 876254528;
assign addr[2547]= 805879757;
assign addr[2548]= 734482665;
assign addr[2549]= 662153826;
assign addr[2550]= 588984994;
assign addr[2551]= 515068990;
assign addr[2552]= 440499581;
assign addr[2553]= 365371365;
assign addr[2554]= 289779648;
assign addr[2555]= 213820322;
assign addr[2556]= 137589750;
assign addr[2557]= 61184634;
assign addr[2558]= -15298099;
assign addr[2559]= -91761426;
assign addr[2560]= -168108346;
assign addr[2561]= -244242007;
assign addr[2562]= -320065829;
assign addr[2563]= -395483624;
assign addr[2564]= -470399716;
assign addr[2565]= -544719071;
assign addr[2566]= -618347408;
assign addr[2567]= -691191324;
assign addr[2568]= -763158411;
assign addr[2569]= -834157373;
assign addr[2570]= -904098143;
assign addr[2571]= -972891995;
assign addr[2572]= -1040451659;
assign addr[2573]= -1106691431;
assign addr[2574]= -1171527280;
assign addr[2575]= -1234876957;
assign addr[2576]= -1296660098;
assign addr[2577]= -1356798326;
assign addr[2578]= -1415215352;
assign addr[2579]= -1471837070;
assign addr[2580]= -1526591649;
assign addr[2581]= -1579409630;
assign addr[2582]= -1630224009;
assign addr[2583]= -1678970324;
assign addr[2584]= -1725586737;
assign addr[2585]= -1770014111;
assign addr[2586]= -1812196087;
assign addr[2587]= -1852079154;
assign addr[2588]= -1889612716;
assign addr[2589]= -1924749160;
assign addr[2590]= -1957443913;
assign addr[2591]= -1987655498;
assign addr[2592]= -2015345591;
assign addr[2593]= -2040479063;
assign addr[2594]= -2063024031;
assign addr[2595]= -2082951896;
assign addr[2596]= -2100237377;
assign addr[2597]= -2114858546;
assign addr[2598]= -2126796855;
assign addr[2599]= -2136037160;
assign addr[2600]= -2142567738;
assign addr[2601]= -2146380306;
assign addr[2602]= -2147470025;
assign addr[2603]= -2145835515;
assign addr[2604]= -2141478848;
assign addr[2605]= -2134405552;
assign addr[2606]= -2124624598;
assign addr[2607]= -2112148396;
assign addr[2608]= -2096992772;
assign addr[2609]= -2079176953;
assign addr[2610]= -2058723538;
assign addr[2611]= -2035658475;
assign addr[2612]= -2010011024;
assign addr[2613]= -1981813720;
assign addr[2614]= -1951102334;
assign addr[2615]= -1917915825;
assign addr[2616]= -1882296293;
assign addr[2617]= -1844288924;
assign addr[2618]= -1803941934;
assign addr[2619]= -1761306505;
assign addr[2620]= -1716436725;
assign addr[2621]= -1669389513;
assign addr[2622]= -1620224553;
assign addr[2623]= -1569004214;
assign addr[2624]= -1515793473;
assign addr[2625]= -1460659832;
assign addr[2626]= -1403673233;
assign addr[2627]= -1344905966;
assign addr[2628]= -1284432584;
assign addr[2629]= -1222329801;
assign addr[2630]= -1158676398;
assign addr[2631]= -1093553126;
assign addr[2632]= -1027042599;
assign addr[2633]= -959229189;
assign addr[2634]= -890198924;
assign addr[2635]= -820039373;
assign addr[2636]= -748839539;
assign addr[2637]= -676689746;
assign addr[2638]= -603681519;
assign addr[2639]= -529907477;
assign addr[2640]= -455461206;
assign addr[2641]= -380437148;
assign addr[2642]= -304930476;
assign addr[2643]= -229036977;
assign addr[2644]= -152852926;
assign addr[2645]= -76474970;
assign addr[2646]= 0;
assign addr[2647]= 76474970;
assign addr[2648]= 152852926;
assign addr[2649]= 229036977;
assign addr[2650]= 304930476;
assign addr[2651]= 380437148;
assign addr[2652]= 455461206;
assign addr[2653]= 529907477;
assign addr[2654]= 603681519;
assign addr[2655]= 676689746;
assign addr[2656]= 748839539;
assign addr[2657]= 820039373;
assign addr[2658]= 890198924;
assign addr[2659]= 959229189;
assign addr[2660]= 1027042599;
assign addr[2661]= 1093553126;
assign addr[2662]= 1158676398;
assign addr[2663]= 1222329801;
assign addr[2664]= 1284432584;
assign addr[2665]= 1344905966;
assign addr[2666]= 1403673233;
assign addr[2667]= 1460659832;
assign addr[2668]= 1515793473;
assign addr[2669]= 1569004214;
assign addr[2670]= 1620224553;
assign addr[2671]= 1669389513;
assign addr[2672]= 1716436725;
assign addr[2673]= 1761306505;
assign addr[2674]= 1803941934;
assign addr[2675]= 1844288924;
assign addr[2676]= 1882296293;
assign addr[2677]= 1917915825;
assign addr[2678]= 1951102334;
assign addr[2679]= 1981813720;
assign addr[2680]= 2010011024;
assign addr[2681]= 2035658475;
assign addr[2682]= 2058723538;
assign addr[2683]= 2079176953;
assign addr[2684]= 2096992772;
assign addr[2685]= 2112148396;
assign addr[2686]= 2124624598;
assign addr[2687]= 2134405552;
assign addr[2688]= 2141478848;
assign addr[2689]= 2145835515;
assign addr[2690]= 2147470025;
assign addr[2691]= 2146380306;
assign addr[2692]= 2142567738;
assign addr[2693]= 2136037160;
assign addr[2694]= 2126796855;
assign addr[2695]= 2114858546;
assign addr[2696]= 2100237377;
assign addr[2697]= 2082951896;
assign addr[2698]= 2063024031;
assign addr[2699]= 2040479063;
assign addr[2700]= 2015345591;
assign addr[2701]= 1987655498;
assign addr[2702]= 1957443913;
assign addr[2703]= 1924749160;
assign addr[2704]= 1889612716;
assign addr[2705]= 1852079154;
assign addr[2706]= 1812196087;
assign addr[2707]= 1770014111;
assign addr[2708]= 1725586737;
assign addr[2709]= 1678970324;
assign addr[2710]= 1630224009;
assign addr[2711]= 1579409630;
assign addr[2712]= 1526591649;
assign addr[2713]= 1471837070;
assign addr[2714]= 1415215352;
assign addr[2715]= 1356798326;
assign addr[2716]= 1296660098;
assign addr[2717]= 1234876957;
assign addr[2718]= 1171527280;
assign addr[2719]= 1106691431;
assign addr[2720]= 1040451659;
assign addr[2721]= 972891995;
assign addr[2722]= 904098143;
assign addr[2723]= 834157373;
assign addr[2724]= 763158411;
assign addr[2725]= 691191324;
assign addr[2726]= 618347408;
assign addr[2727]= 544719071;
assign addr[2728]= 470399716;
assign addr[2729]= 395483624;
assign addr[2730]= 320065829;
assign addr[2731]= 244242007;
assign addr[2732]= 168108346;
assign addr[2733]= 91761426;
assign addr[2734]= 15298099;
assign addr[2735]= -61184634;
assign addr[2736]= -137589750;
assign addr[2737]= -213820322;
assign addr[2738]= -289779648;
assign addr[2739]= -365371365;
assign addr[2740]= -440499581;
assign addr[2741]= -515068990;
assign addr[2742]= -588984994;
assign addr[2743]= -662153826;
assign addr[2744]= -734482665;
assign addr[2745]= -805879757;
assign addr[2746]= -876254528;
assign addr[2747]= -945517704;
assign addr[2748]= -1013581418;
assign addr[2749]= -1080359326;
assign addr[2750]= -1145766716;
assign addr[2751]= -1209720613;
assign addr[2752]= -1272139887;
assign addr[2753]= -1332945355;
assign addr[2754]= -1392059879;
assign addr[2755]= -1449408469;
assign addr[2756]= -1504918373;
assign addr[2757]= -1558519173;
assign addr[2758]= -1610142873;
assign addr[2759]= -1659723983;
assign addr[2760]= -1707199606;
assign addr[2761]= -1752509516;
assign addr[2762]= -1795596234;
assign addr[2763]= -1836405100;
assign addr[2764]= -1874884346;
assign addr[2765]= -1910985158;
assign addr[2766]= -1944661739;
assign addr[2767]= -1975871368;
assign addr[2768]= -2004574453;
assign addr[2769]= -2030734582;
assign addr[2770]= -2054318569;
assign addr[2771]= -2075296495;
assign addr[2772]= -2093641749;
assign addr[2773]= -2109331059;
assign addr[2774]= -2122344521;
assign addr[2775]= -2132665626;
assign addr[2776]= -2140281282;
assign addr[2777]= -2145181827;
assign addr[2778]= -2147361045;
assign addr[2779]= -2146816171;
assign addr[2780]= -2143547897;
assign addr[2781]= -2137560369;
assign addr[2782]= -2128861181;
assign addr[2783]= -2117461370;
assign addr[2784]= -2103375398;
assign addr[2785]= -2086621133;
assign addr[2786]= -2067219829;
assign addr[2787]= -2045196100;
assign addr[2788]= -2020577882;
assign addr[2789]= -1993396407;
assign addr[2790]= -1963686155;
assign addr[2791]= -1931484818;
assign addr[2792]= -1896833245;
assign addr[2793]= -1859775393;
assign addr[2794]= -1820358275;
assign addr[2795]= -1778631892;
assign addr[2796]= -1734649179;
assign addr[2797]= -1688465931;
assign addr[2798]= -1640140734;
assign addr[2799]= -1589734894;
assign addr[2800]= -1537312353;
assign addr[2801]= -1482939614;
assign addr[2802]= -1426685652;
assign addr[2803]= -1368621831;
assign addr[2804]= -1308821808;
assign addr[2805]= -1247361445;
assign addr[2806]= -1184318708;
assign addr[2807]= -1119773573;
assign addr[2808]= -1053807919;
assign addr[2809]= -986505429;
assign addr[2810]= -917951481;
assign addr[2811]= -848233042;
assign addr[2812]= -777438554;
assign addr[2813]= -705657826;
assign addr[2814]= -632981917;
assign addr[2815]= -559503022;
assign addr[2816]= -485314355;
assign addr[2817]= -410510029;
assign addr[2818]= -335184940;
assign addr[2819]= -259434643;
assign addr[2820]= -183355234;
assign addr[2821]= -107043224;
assign addr[2822]= -30595422;
assign addr[2823]= 45891193;
assign addr[2824]= 122319591;
assign addr[2825]= 198592817;
assign addr[2826]= 274614114;
assign addr[2827]= 350287041;
assign addr[2828]= 425515602;
assign addr[2829]= 500204365;
assign addr[2830]= 574258580;
assign addr[2831]= 647584304;
assign addr[2832]= 720088517;
assign addr[2833]= 791679244;
assign addr[2834]= 862265664;
assign addr[2835]= 931758235;
assign addr[2836]= 1000068799;
assign addr[2837]= 1067110699;
assign addr[2838]= 1132798888;
assign addr[2839]= 1197050035;
assign addr[2840]= 1259782632;
assign addr[2841]= 1320917099;
assign addr[2842]= 1380375881;
assign addr[2843]= 1438083551;
assign addr[2844]= 1493966902;
assign addr[2845]= 1547955041;
assign addr[2846]= 1599979481;
assign addr[2847]= 1649974225;
assign addr[2848]= 1697875851;
assign addr[2849]= 1743623590;
assign addr[2850]= 1787159411;
assign addr[2851]= 1828428082;
assign addr[2852]= 1867377253;
assign addr[2853]= 1903957513;
assign addr[2854]= 1938122457;
assign addr[2855]= 1969828744;
assign addr[2856]= 1999036154;
assign addr[2857]= 2025707632;
assign addr[2858]= 2049809346;
assign addr[2859]= 2071310720;
assign addr[2860]= 2090184478;
assign addr[2861]= 2106406677;
assign addr[2862]= 2119956737;
assign addr[2863]= 2130817471;
assign addr[2864]= 2138975100;
assign addr[2865]= 2144419275;
assign addr[2866]= 2147143090;
assign addr[2867]= 2147143090;
assign addr[2868]= 2144419275;
assign addr[2869]= 2138975100;
assign addr[2870]= 2130817471;
assign addr[2871]= 2119956737;
assign addr[2872]= 2106406677;
assign addr[2873]= 2090184478;
assign addr[2874]= 2071310720;
assign addr[2875]= 2049809346;
assign addr[2876]= 2025707632;
assign addr[2877]= 1999036154;
assign addr[2878]= 1969828744;
assign addr[2879]= 1938122457;
assign addr[2880]= 1903957513;
assign addr[2881]= 1867377253;
assign addr[2882]= 1828428082;
assign addr[2883]= 1787159411;
assign addr[2884]= 1743623590;
assign addr[2885]= 1697875851;
assign addr[2886]= 1649974225;
assign addr[2887]= 1599979481;
assign addr[2888]= 1547955041;
assign addr[2889]= 1493966902;
assign addr[2890]= 1438083551;
assign addr[2891]= 1380375881;
assign addr[2892]= 1320917099;
assign addr[2893]= 1259782632;
assign addr[2894]= 1197050035;
assign addr[2895]= 1132798888;
assign addr[2896]= 1067110699;
assign addr[2897]= 1000068799;
assign addr[2898]= 931758235;
assign addr[2899]= 862265664;
assign addr[2900]= 791679244;
assign addr[2901]= 720088517;
assign addr[2902]= 647584304;
assign addr[2903]= 574258580;
assign addr[2904]= 500204365;
assign addr[2905]= 425515602;
assign addr[2906]= 350287041;
assign addr[2907]= 274614114;
assign addr[2908]= 198592817;
assign addr[2909]= 122319591;
assign addr[2910]= 45891193;
assign addr[2911]= -30595422;
assign addr[2912]= -107043224;
assign addr[2913]= -183355234;
assign addr[2914]= -259434643;
assign addr[2915]= -335184940;
assign addr[2916]= -410510029;
assign addr[2917]= -485314355;
assign addr[2918]= -559503022;
assign addr[2919]= -632981917;
assign addr[2920]= -705657826;
assign addr[2921]= -777438554;
assign addr[2922]= -848233042;
assign addr[2923]= -917951481;
assign addr[2924]= -986505429;
assign addr[2925]= -1053807919;
assign addr[2926]= -1119773573;
assign addr[2927]= -1184318708;
assign addr[2928]= -1247361445;
assign addr[2929]= -1308821808;
assign addr[2930]= -1368621831;
assign addr[2931]= -1426685652;
assign addr[2932]= -1482939614;
assign addr[2933]= -1537312353;
assign addr[2934]= -1589734894;
assign addr[2935]= -1640140734;
assign addr[2936]= -1688465931;
assign addr[2937]= -1734649179;
assign addr[2938]= -1778631892;
assign addr[2939]= -1820358275;
assign addr[2940]= -1859775393;
assign addr[2941]= -1896833245;
assign addr[2942]= -1931484818;
assign addr[2943]= -1963686155;
assign addr[2944]= -1993396407;
assign addr[2945]= -2020577882;
assign addr[2946]= -2045196100;
assign addr[2947]= -2067219829;
assign addr[2948]= -2086621133;
assign addr[2949]= -2103375398;
assign addr[2950]= -2117461370;
assign addr[2951]= -2128861181;
assign addr[2952]= -2137560369;
assign addr[2953]= -2143547897;
assign addr[2954]= -2146816171;
assign addr[2955]= -2147361045;
assign addr[2956]= -2145181827;
assign addr[2957]= -2140281282;
assign addr[2958]= -2132665626;
assign addr[2959]= -2122344521;
assign addr[2960]= -2109331059;
assign addr[2961]= -2093641749;
assign addr[2962]= -2075296495;
assign addr[2963]= -2054318569;
assign addr[2964]= -2030734582;
assign addr[2965]= -2004574453;
assign addr[2966]= -1975871368;
assign addr[2967]= -1944661739;
assign addr[2968]= -1910985158;
assign addr[2969]= -1874884346;
assign addr[2970]= -1836405100;
assign addr[2971]= -1795596234;
assign addr[2972]= -1752509516;
assign addr[2973]= -1707199606;
assign addr[2974]= -1659723983;
assign addr[2975]= -1610142873;
assign addr[2976]= -1558519173;
assign addr[2977]= -1504918373;
assign addr[2978]= -1449408469;
assign addr[2979]= -1392059879;
assign addr[2980]= -1332945355;
assign addr[2981]= -1272139887;
assign addr[2982]= -1209720613;
assign addr[2983]= -1145766716;
assign addr[2984]= -1080359326;
assign addr[2985]= -1013581418;
assign addr[2986]= -945517704;
assign addr[2987]= -876254528;
assign addr[2988]= -805879757;
assign addr[2989]= -734482665;
assign addr[2990]= -662153826;
assign addr[2991]= -588984994;
assign addr[2992]= -515068990;
assign addr[2993]= -440499581;
assign addr[2994]= -365371365;
assign addr[2995]= -289779648;
assign addr[2996]= -213820322;
assign addr[2997]= -137589750;
assign addr[2998]= -61184634;
assign addr[2999]= 15298099;
assign addr[3000]= 91761426;
assign addr[3001]= 168108346;
assign addr[3002]= 244242007;
assign addr[3003]= 320065829;
assign addr[3004]= 395483624;
assign addr[3005]= 470399716;
assign addr[3006]= 544719071;
assign addr[3007]= 618347408;
assign addr[3008]= 691191324;
assign addr[3009]= 763158411;
assign addr[3010]= 834157373;
assign addr[3011]= 904098143;
assign addr[3012]= 972891995;
assign addr[3013]= 1040451659;
assign addr[3014]= 1106691431;
assign addr[3015]= 1171527280;
assign addr[3016]= 1234876957;
assign addr[3017]= 1296660098;
assign addr[3018]= 1356798326;
assign addr[3019]= 1415215352;
assign addr[3020]= 1471837070;
assign addr[3021]= 1526591649;
assign addr[3022]= 1579409630;
assign addr[3023]= 1630224009;
assign addr[3024]= 1678970324;
assign addr[3025]= 1725586737;
assign addr[3026]= 1770014111;
assign addr[3027]= 1812196087;
assign addr[3028]= 1852079154;
assign addr[3029]= 1889612716;
assign addr[3030]= 1924749160;
assign addr[3031]= 1957443913;
assign addr[3032]= 1987655498;
assign addr[3033]= 2015345591;
assign addr[3034]= 2040479063;
assign addr[3035]= 2063024031;
assign addr[3036]= 2082951896;
assign addr[3037]= 2100237377;
assign addr[3038]= 2114858546;
assign addr[3039]= 2126796855;
assign addr[3040]= 2136037160;
assign addr[3041]= 2142567738;
assign addr[3042]= 2146380306;
assign addr[3043]= 2147470025;
assign addr[3044]= 2145835515;
assign addr[3045]= 2141478848;
assign addr[3046]= 2134405552;
assign addr[3047]= 2124624598;
assign addr[3048]= 2112148396;
assign addr[3049]= 2096992772;
assign addr[3050]= 2079176953;
assign addr[3051]= 2058723538;
assign addr[3052]= 2035658475;
assign addr[3053]= 2010011024;
assign addr[3054]= 1981813720;
assign addr[3055]= 1951102334;
assign addr[3056]= 1917915825;
assign addr[3057]= 1882296293;
assign addr[3058]= 1844288924;
assign addr[3059]= 1803941934;
assign addr[3060]= 1761306505;
assign addr[3061]= 1716436725;
assign addr[3062]= 1669389513;
assign addr[3063]= 1620224553;
assign addr[3064]= 1569004214;
assign addr[3065]= 1515793473;
assign addr[3066]= 1460659832;
assign addr[3067]= 1403673233;
assign addr[3068]= 1344905966;
assign addr[3069]= 1284432584;
assign addr[3070]= 1222329801;
assign addr[3071]= 1158676398;
assign addr[3072]= 1093553126;
assign addr[3073]= 1027042599;
assign addr[3074]= 959229189;
assign addr[3075]= 890198924;
assign addr[3076]= 820039373;
assign addr[3077]= 748839539;
assign addr[3078]= 676689746;
assign addr[3079]= 603681519;
assign addr[3080]= 529907477;
assign addr[3081]= 455461206;
assign addr[3082]= 380437148;
assign addr[3083]= 304930476;
assign addr[3084]= 229036977;
assign addr[3085]= 152852926;
assign addr[3086]= 76474970;
assign addr[3087]= 0;
assign addr[3088]= -76474970;
assign addr[3089]= -152852926;
assign addr[3090]= -229036977;
assign addr[3091]= -304930476;
assign addr[3092]= -380437148;
assign addr[3093]= -455461206;
assign addr[3094]= -529907477;
assign addr[3095]= -603681519;
assign addr[3096]= -676689746;
assign addr[3097]= -748839539;
assign addr[3098]= -820039373;
assign addr[3099]= -890198924;
assign addr[3100]= -959229189;
assign addr[3101]= -1027042599;
assign addr[3102]= -1093553126;
assign addr[3103]= -1158676398;
assign addr[3104]= -1222329801;
assign addr[3105]= -1284432584;
assign addr[3106]= -1344905966;
assign addr[3107]= -1403673233;
assign addr[3108]= -1460659832;
assign addr[3109]= -1515793473;
assign addr[3110]= -1569004214;
assign addr[3111]= -1620224553;
assign addr[3112]= -1669389513;
assign addr[3113]= -1716436725;
assign addr[3114]= -1761306505;
assign addr[3115]= -1803941934;
assign addr[3116]= -1844288924;
assign addr[3117]= -1882296293;
assign addr[3118]= -1917915825;
assign addr[3119]= -1951102334;
assign addr[3120]= -1981813720;
assign addr[3121]= -2010011024;
assign addr[3122]= -2035658475;
assign addr[3123]= -2058723538;
assign addr[3124]= -2079176953;
assign addr[3125]= -2096992772;
assign addr[3126]= -2112148396;
assign addr[3127]= -2124624598;
assign addr[3128]= -2134405552;
assign addr[3129]= -2141478848;
assign addr[3130]= -2145835515;
assign addr[3131]= -2147470025;
assign addr[3132]= -2146380306;
assign addr[3133]= -2142567738;
assign addr[3134]= -2136037160;
assign addr[3135]= -2126796855;
assign addr[3136]= -2114858546;
assign addr[3137]= -2100237377;
assign addr[3138]= -2082951896;
assign addr[3139]= -2063024031;
assign addr[3140]= -2040479063;
assign addr[3141]= -2015345591;
assign addr[3142]= -1987655498;
assign addr[3143]= -1957443913;
assign addr[3144]= -1924749160;
assign addr[3145]= -1889612716;
assign addr[3146]= -1852079154;
assign addr[3147]= -1812196087;
assign addr[3148]= -1770014111;
assign addr[3149]= -1725586737;
assign addr[3150]= -1678970324;
assign addr[3151]= -1630224009;
assign addr[3152]= -1579409630;
assign addr[3153]= -1526591649;
assign addr[3154]= -1471837070;
assign addr[3155]= -1415215352;
assign addr[3156]= -1356798326;
assign addr[3157]= -1296660098;
assign addr[3158]= -1234876957;
assign addr[3159]= -1171527280;
assign addr[3160]= -1106691431;
assign addr[3161]= -1040451659;
assign addr[3162]= -972891995;
assign addr[3163]= -904098143;
assign addr[3164]= -834157373;
assign addr[3165]= -763158411;
assign addr[3166]= -691191324;
assign addr[3167]= -618347408;
assign addr[3168]= -544719071;
assign addr[3169]= -470399716;
assign addr[3170]= -395483624;
assign addr[3171]= -320065829;
assign addr[3172]= -244242007;
assign addr[3173]= -168108346;
assign addr[3174]= -91761426;
assign addr[3175]= -15298099;
assign addr[3176]= 61184634;
assign addr[3177]= 137589750;
assign addr[3178]= 213820322;
assign addr[3179]= 289779648;
assign addr[3180]= 365371365;
assign addr[3181]= 440499581;
assign addr[3182]= 515068990;
assign addr[3183]= 588984994;
assign addr[3184]= 662153826;
assign addr[3185]= 734482665;
assign addr[3186]= 805879757;
assign addr[3187]= 876254528;
assign addr[3188]= 945517704;
assign addr[3189]= 1013581418;
assign addr[3190]= 1080359326;
assign addr[3191]= 1145766716;
assign addr[3192]= 1209720613;
assign addr[3193]= 1272139887;
assign addr[3194]= 1332945355;
assign addr[3195]= 1392059879;
assign addr[3196]= 1449408469;
assign addr[3197]= 1504918373;
assign addr[3198]= 1558519173;
assign addr[3199]= 1610142873;
assign addr[3200]= 1659723983;
assign addr[3201]= 1707199606;
assign addr[3202]= 1752509516;
assign addr[3203]= 1795596234;
assign addr[3204]= 1836405100;
assign addr[3205]= 1874884346;
assign addr[3206]= 1910985158;
assign addr[3207]= 1944661739;
assign addr[3208]= 1975871368;
assign addr[3209]= 2004574453;
assign addr[3210]= 2030734582;
assign addr[3211]= 2054318569;
assign addr[3212]= 2075296495;
assign addr[3213]= 2093641749;
assign addr[3214]= 2109331059;
assign addr[3215]= 2122344521;
assign addr[3216]= 2132665626;
assign addr[3217]= 2140281282;
assign addr[3218]= 2145181827;
assign addr[3219]= 2147361045;
assign addr[3220]= 2146816171;
assign addr[3221]= 2143547897;
assign addr[3222]= 2137560369;
assign addr[3223]= 2128861181;
assign addr[3224]= 2117461370;
assign addr[3225]= 2103375398;
assign addr[3226]= 2086621133;
assign addr[3227]= 2067219829;
assign addr[3228]= 2045196100;
assign addr[3229]= 2020577882;
assign addr[3230]= 1993396407;
assign addr[3231]= 1963686155;
assign addr[3232]= 1931484818;
assign addr[3233]= 1896833245;
assign addr[3234]= 1859775393;
assign addr[3235]= 1820358275;
assign addr[3236]= 1778631892;
assign addr[3237]= 1734649179;
assign addr[3238]= 1688465931;
assign addr[3239]= 1640140734;
assign addr[3240]= 1589734894;
assign addr[3241]= 1537312353;
assign addr[3242]= 1482939614;
assign addr[3243]= 1426685652;
assign addr[3244]= 1368621831;
assign addr[3245]= 1308821808;
assign addr[3246]= 1247361445;
assign addr[3247]= 1184318708;
assign addr[3248]= 1119773573;
assign addr[3249]= 1053807919;
assign addr[3250]= 986505429;
assign addr[3251]= 917951481;
assign addr[3252]= 848233042;
assign addr[3253]= 777438554;
assign addr[3254]= 705657826;
assign addr[3255]= 632981917;
assign addr[3256]= 559503022;
assign addr[3257]= 485314355;
assign addr[3258]= 410510029;
assign addr[3259]= 335184940;
assign addr[3260]= 259434643;
assign addr[3261]= 183355234;
assign addr[3262]= 107043224;
assign addr[3263]= 30595422;
assign addr[3264]= -45891193;
assign addr[3265]= -122319591;
assign addr[3266]= -198592817;
assign addr[3267]= -274614114;
assign addr[3268]= -350287041;
assign addr[3269]= -425515602;
assign addr[3270]= -500204365;
assign addr[3271]= -574258580;
assign addr[3272]= -647584304;
assign addr[3273]= -720088517;
assign addr[3274]= -791679244;
assign addr[3275]= -862265664;
assign addr[3276]= -931758235;
assign addr[3277]= -1000068799;
assign addr[3278]= -1067110699;
assign addr[3279]= -1132798888;
assign addr[3280]= -1197050035;
assign addr[3281]= -1259782632;
assign addr[3282]= -1320917099;
assign addr[3283]= -1380375881;
assign addr[3284]= -1438083551;
assign addr[3285]= -1493966902;
assign addr[3286]= -1547955041;
assign addr[3287]= -1599979481;
assign addr[3288]= -1649974225;
assign addr[3289]= -1697875851;
assign addr[3290]= -1743623590;
assign addr[3291]= -1787159411;
assign addr[3292]= -1828428082;
assign addr[3293]= -1867377253;
assign addr[3294]= -1903957513;
assign addr[3295]= -1938122457;
assign addr[3296]= -1969828744;
assign addr[3297]= -1999036154;
assign addr[3298]= -2025707632;
assign addr[3299]= -2049809346;
assign addr[3300]= -2071310720;
assign addr[3301]= -2090184478;
assign addr[3302]= -2106406677;
assign addr[3303]= -2119956737;
assign addr[3304]= -2130817471;
assign addr[3305]= -2138975100;
assign addr[3306]= -2144419275;
assign addr[3307]= -2147143090;
assign addr[3308]= -2147143090;
assign addr[3309]= -2144419275;
assign addr[3310]= -2138975100;
assign addr[3311]= -2130817471;
assign addr[3312]= -2119956737;
assign addr[3313]= -2106406677;
assign addr[3314]= -2090184478;
assign addr[3315]= -2071310720;
assign addr[3316]= -2049809346;
assign addr[3317]= -2025707632;
assign addr[3318]= -1999036154;
assign addr[3319]= -1969828744;
assign addr[3320]= -1938122457;
assign addr[3321]= -1903957513;
assign addr[3322]= -1867377253;
assign addr[3323]= -1828428082;
assign addr[3324]= -1787159411;
assign addr[3325]= -1743623590;
assign addr[3326]= -1697875851;
assign addr[3327]= -1649974225;
assign addr[3328]= -1599979481;
assign addr[3329]= -1547955041;
assign addr[3330]= -1493966902;
assign addr[3331]= -1438083551;
assign addr[3332]= -1380375881;
assign addr[3333]= -1320917099;
assign addr[3334]= -1259782632;
assign addr[3335]= -1197050035;
assign addr[3336]= -1132798888;
assign addr[3337]= -1067110699;
assign addr[3338]= -1000068799;
assign addr[3339]= -931758235;
assign addr[3340]= -862265664;
assign addr[3341]= -791679244;
assign addr[3342]= -720088517;
assign addr[3343]= -647584304;
assign addr[3344]= -574258580;
assign addr[3345]= -500204365;
assign addr[3346]= -425515602;
assign addr[3347]= -350287041;
assign addr[3348]= -274614114;
assign addr[3349]= -198592817;
assign addr[3350]= -122319591;
assign addr[3351]= -45891193;
assign addr[3352]= 30595422;
assign addr[3353]= 107043224;
assign addr[3354]= 183355234;
assign addr[3355]= 259434643;
assign addr[3356]= 335184940;
assign addr[3357]= 410510029;
assign addr[3358]= 485314355;
assign addr[3359]= 559503022;
assign addr[3360]= 632981917;
assign addr[3361]= 705657826;
assign addr[3362]= 777438554;
assign addr[3363]= 848233042;
assign addr[3364]= 917951481;
assign addr[3365]= 986505429;
assign addr[3366]= 1053807919;
assign addr[3367]= 1119773573;
assign addr[3368]= 1184318708;
assign addr[3369]= 1247361445;
assign addr[3370]= 1308821808;
assign addr[3371]= 1368621831;
assign addr[3372]= 1426685652;
assign addr[3373]= 1482939614;
assign addr[3374]= 1537312353;
assign addr[3375]= 1589734894;
assign addr[3376]= 1640140734;
assign addr[3377]= 1688465931;
assign addr[3378]= 1734649179;
assign addr[3379]= 1778631892;
assign addr[3380]= 1820358275;
assign addr[3381]= 1859775393;
assign addr[3382]= 1896833245;
assign addr[3383]= 1931484818;
assign addr[3384]= 1963686155;
assign addr[3385]= 1993396407;
assign addr[3386]= 2020577882;
assign addr[3387]= 2045196100;
assign addr[3388]= 2067219829;
assign addr[3389]= 2086621133;
assign addr[3390]= 2103375398;
assign addr[3391]= 2117461370;
assign addr[3392]= 2128861181;
assign addr[3393]= 2137560369;
assign addr[3394]= 2143547897;
assign addr[3395]= 2146816171;
assign addr[3396]= 2147361045;
assign addr[3397]= 2145181827;
assign addr[3398]= 2140281282;
assign addr[3399]= 2132665626;
assign addr[3400]= 2122344521;
assign addr[3401]= 2109331059;
assign addr[3402]= 2093641749;
assign addr[3403]= 2075296495;
assign addr[3404]= 2054318569;
assign addr[3405]= 2030734582;
assign addr[3406]= 2004574453;
assign addr[3407]= 1975871368;
assign addr[3408]= 1944661739;
assign addr[3409]= 1910985158;
assign addr[3410]= 1874884346;
assign addr[3411]= 1836405100;
assign addr[3412]= 1795596234;
assign addr[3413]= 1752509516;
assign addr[3414]= 1707199606;
assign addr[3415]= 1659723983;
assign addr[3416]= 1610142873;
assign addr[3417]= 1558519173;
assign addr[3418]= 1504918373;
assign addr[3419]= 1449408469;
assign addr[3420]= 1392059879;
assign addr[3421]= 1332945355;
assign addr[3422]= 1272139887;
assign addr[3423]= 1209720613;
assign addr[3424]= 1145766716;
assign addr[3425]= 1080359326;
assign addr[3426]= 1013581418;
assign addr[3427]= 945517704;
assign addr[3428]= 876254528;
assign addr[3429]= 805879757;
assign addr[3430]= 734482665;
assign addr[3431]= 662153826;
assign addr[3432]= 588984994;
assign addr[3433]= 515068990;
assign addr[3434]= 440499581;
assign addr[3435]= 365371365;
assign addr[3436]= 289779648;
assign addr[3437]= 213820322;
assign addr[3438]= 137589750;
assign addr[3439]= 61184634;
assign addr[3440]= -15298099;
assign addr[3441]= -91761426;
assign addr[3442]= -168108346;
assign addr[3443]= -244242007;
assign addr[3444]= -320065829;
assign addr[3445]= -395483624;
assign addr[3446]= -470399716;
assign addr[3447]= -544719071;
assign addr[3448]= -618347408;
assign addr[3449]= -691191324;
assign addr[3450]= -763158411;
assign addr[3451]= -834157373;
assign addr[3452]= -904098143;
assign addr[3453]= -972891995;
assign addr[3454]= -1040451659;
assign addr[3455]= -1106691431;
assign addr[3456]= -1171527280;
assign addr[3457]= -1234876957;
assign addr[3458]= -1296660098;
assign addr[3459]= -1356798326;
assign addr[3460]= -1415215352;
assign addr[3461]= -1471837070;
assign addr[3462]= -1526591649;
assign addr[3463]= -1579409630;
assign addr[3464]= -1630224009;
assign addr[3465]= -1678970324;
assign addr[3466]= -1725586737;
assign addr[3467]= -1770014111;
assign addr[3468]= -1812196087;
assign addr[3469]= -1852079154;
assign addr[3470]= -1889612716;
assign addr[3471]= -1924749160;
assign addr[3472]= -1957443913;
assign addr[3473]= -1987655498;
assign addr[3474]= -2015345591;
assign addr[3475]= -2040479063;
assign addr[3476]= -2063024031;
assign addr[3477]= -2082951896;
assign addr[3478]= -2100237377;
assign addr[3479]= -2114858546;
assign addr[3480]= -2126796855;
assign addr[3481]= -2136037160;
assign addr[3482]= -2142567738;
assign addr[3483]= -2146380306;
assign addr[3484]= -2147470025;
assign addr[3485]= -2145835515;
assign addr[3486]= -2141478848;
assign addr[3487]= -2134405552;
assign addr[3488]= -2124624598;
assign addr[3489]= -2112148396;
assign addr[3490]= -2096992772;
assign addr[3491]= -2079176953;
assign addr[3492]= -2058723538;
assign addr[3493]= -2035658475;
assign addr[3494]= -2010011024;
assign addr[3495]= -1981813720;
assign addr[3496]= -1951102334;
assign addr[3497]= -1917915825;
assign addr[3498]= -1882296293;
assign addr[3499]= -1844288924;
assign addr[3500]= -1803941934;
assign addr[3501]= -1761306505;
assign addr[3502]= -1716436725;
assign addr[3503]= -1669389513;
assign addr[3504]= -1620224553;
assign addr[3505]= -1569004214;
assign addr[3506]= -1515793473;
assign addr[3507]= -1460659832;
assign addr[3508]= -1403673233;
assign addr[3509]= -1344905966;
assign addr[3510]= -1284432584;
assign addr[3511]= -1222329801;
assign addr[3512]= -1158676398;
assign addr[3513]= -1093553126;
assign addr[3514]= -1027042599;
assign addr[3515]= -959229189;
assign addr[3516]= -890198924;
assign addr[3517]= -820039373;
assign addr[3518]= -748839539;
assign addr[3519]= -676689746;
assign addr[3520]= -603681519;
assign addr[3521]= -529907477;
assign addr[3522]= -455461206;
assign addr[3523]= -380437148;
assign addr[3524]= -304930476;
assign addr[3525]= -229036977;
assign addr[3526]= -152852926;
assign addr[3527]= -76474970;
assign addr[3528]= 0;
assign addr[3529]= 76474970;
assign addr[3530]= 152852926;
assign addr[3531]= 229036977;
assign addr[3532]= 304930476;
assign addr[3533]= 380437148;
assign addr[3534]= 455461206;
assign addr[3535]= 529907477;
assign addr[3536]= 603681519;
assign addr[3537]= 676689746;
assign addr[3538]= 748839539;
assign addr[3539]= 820039373;
assign addr[3540]= 890198924;
assign addr[3541]= 959229189;
assign addr[3542]= 1027042599;
assign addr[3543]= 1093553126;
assign addr[3544]= 1158676398;
assign addr[3545]= 1222329801;
assign addr[3546]= 1284432584;
assign addr[3547]= 1344905966;
assign addr[3548]= 1403673233;
assign addr[3549]= 1460659832;
assign addr[3550]= 1515793473;
assign addr[3551]= 1569004214;
assign addr[3552]= 1620224553;
assign addr[3553]= 1669389513;
assign addr[3554]= 1716436725;
assign addr[3555]= 1761306505;
assign addr[3556]= 1803941934;
assign addr[3557]= 1844288924;
assign addr[3558]= 1882296293;
assign addr[3559]= 1917915825;
assign addr[3560]= 1951102334;
assign addr[3561]= 1981813720;
assign addr[3562]= 2010011024;
assign addr[3563]= 2035658475;
assign addr[3564]= 2058723538;
assign addr[3565]= 2079176953;
assign addr[3566]= 2096992772;
assign addr[3567]= 2112148396;
assign addr[3568]= 2124624598;
assign addr[3569]= 2134405552;
assign addr[3570]= 2141478848;
assign addr[3571]= 2145835515;
assign addr[3572]= 2147470025;
assign addr[3573]= 2146380306;
assign addr[3574]= 2142567738;
assign addr[3575]= 2136037160;
assign addr[3576]= 2126796855;
assign addr[3577]= 2114858546;
assign addr[3578]= 2100237377;
assign addr[3579]= 2082951896;
assign addr[3580]= 2063024031;
assign addr[3581]= 2040479063;
assign addr[3582]= 2015345591;
assign addr[3583]= 1987655498;
assign addr[3584]= 1957443913;
assign addr[3585]= 1924749160;
assign addr[3586]= 1889612716;
assign addr[3587]= 1852079154;
assign addr[3588]= 1812196087;
assign addr[3589]= 1770014111;
assign addr[3590]= 1725586737;
assign addr[3591]= 1678970324;
assign addr[3592]= 1630224009;
assign addr[3593]= 1579409630;
assign addr[3594]= 1526591649;
assign addr[3595]= 1471837070;
assign addr[3596]= 1415215352;
assign addr[3597]= 1356798326;
assign addr[3598]= 1296660098;
assign addr[3599]= 1234876957;
assign addr[3600]= 1171527280;
assign addr[3601]= 1106691431;
assign addr[3602]= 1040451659;
assign addr[3603]= 972891995;
assign addr[3604]= 904098143;
assign addr[3605]= 834157373;
assign addr[3606]= 763158411;
assign addr[3607]= 691191324;
assign addr[3608]= 618347408;
assign addr[3609]= 544719071;
assign addr[3610]= 470399716;
assign addr[3611]= 395483624;
assign addr[3612]= 320065829;
assign addr[3613]= 244242007;
assign addr[3614]= 168108346;
assign addr[3615]= 91761426;
assign addr[3616]= 15298099;
assign addr[3617]= -61184634;
assign addr[3618]= -137589750;
assign addr[3619]= -213820322;
assign addr[3620]= -289779648;
assign addr[3621]= -365371365;
assign addr[3622]= -440499581;
assign addr[3623]= -515068990;
assign addr[3624]= -588984994;
assign addr[3625]= -662153826;
assign addr[3626]= -734482665;
assign addr[3627]= -805879757;
assign addr[3628]= -876254528;
assign addr[3629]= -945517704;
assign addr[3630]= -1013581418;
assign addr[3631]= -1080359326;
assign addr[3632]= -1145766716;
assign addr[3633]= -1209720613;
assign addr[3634]= -1272139887;
assign addr[3635]= -1332945355;
assign addr[3636]= -1392059879;
assign addr[3637]= -1449408469;
assign addr[3638]= -1504918373;
assign addr[3639]= -1558519173;
assign addr[3640]= -1610142873;
assign addr[3641]= -1659723983;
assign addr[3642]= -1707199606;
assign addr[3643]= -1752509516;
assign addr[3644]= -1795596234;
assign addr[3645]= -1836405100;
assign addr[3646]= -1874884346;
assign addr[3647]= -1910985158;
assign addr[3648]= -1944661739;
assign addr[3649]= -1975871368;
assign addr[3650]= -2004574453;
assign addr[3651]= -2030734582;
assign addr[3652]= -2054318569;
assign addr[3653]= -2075296495;
assign addr[3654]= -2093641749;
assign addr[3655]= -2109331059;
assign addr[3656]= -2122344521;
assign addr[3657]= -2132665626;
assign addr[3658]= -2140281282;
assign addr[3659]= -2145181827;
assign addr[3660]= -2147361045;
assign addr[3661]= -2146816171;
assign addr[3662]= -2143547897;
assign addr[3663]= -2137560369;
assign addr[3664]= -2128861181;
assign addr[3665]= -2117461370;
assign addr[3666]= -2103375398;
assign addr[3667]= -2086621133;
assign addr[3668]= -2067219829;
assign addr[3669]= -2045196100;
assign addr[3670]= -2020577882;
assign addr[3671]= -1993396407;
assign addr[3672]= -1963686155;
assign addr[3673]= -1931484818;
assign addr[3674]= -1896833245;
assign addr[3675]= -1859775393;
assign addr[3676]= -1820358275;
assign addr[3677]= -1778631892;
assign addr[3678]= -1734649179;
assign addr[3679]= -1688465931;
assign addr[3680]= -1640140734;
assign addr[3681]= -1589734894;
assign addr[3682]= -1537312353;
assign addr[3683]= -1482939614;
assign addr[3684]= -1426685652;
assign addr[3685]= -1368621831;
assign addr[3686]= -1308821808;
assign addr[3687]= -1247361445;
assign addr[3688]= -1184318708;
assign addr[3689]= -1119773573;
assign addr[3690]= -1053807919;
assign addr[3691]= -986505429;
assign addr[3692]= -917951481;
assign addr[3693]= -848233042;
assign addr[3694]= -777438554;
assign addr[3695]= -705657826;
assign addr[3696]= -632981917;
assign addr[3697]= -559503022;
assign addr[3698]= -485314355;
assign addr[3699]= -410510029;
assign addr[3700]= -335184940;
assign addr[3701]= -259434643;
assign addr[3702]= -183355234;
assign addr[3703]= -107043224;
assign addr[3704]= -30595422;
assign addr[3705]= 45891193;
assign addr[3706]= 122319591;
assign addr[3707]= 198592817;
assign addr[3708]= 274614114;
assign addr[3709]= 350287041;
assign addr[3710]= 425515602;
assign addr[3711]= 500204365;
assign addr[3712]= 574258580;
assign addr[3713]= 647584304;
assign addr[3714]= 720088517;
assign addr[3715]= 791679244;
assign addr[3716]= 862265664;
assign addr[3717]= 931758235;
assign addr[3718]= 1000068799;
assign addr[3719]= 1067110699;
assign addr[3720]= 1132798888;
assign addr[3721]= 1197050035;
assign addr[3722]= 1259782632;
assign addr[3723]= 1320917099;
assign addr[3724]= 1380375881;
assign addr[3725]= 1438083551;
assign addr[3726]= 1493966902;
assign addr[3727]= 1547955041;
assign addr[3728]= 1599979481;
assign addr[3729]= 1649974225;
assign addr[3730]= 1697875851;
assign addr[3731]= 1743623590;
assign addr[3732]= 1787159411;
assign addr[3733]= 1828428082;
assign addr[3734]= 1867377253;
assign addr[3735]= 1903957513;
assign addr[3736]= 1938122457;
assign addr[3737]= 1969828744;
assign addr[3738]= 1999036154;
assign addr[3739]= 2025707632;
assign addr[3740]= 2049809346;
assign addr[3741]= 2071310720;
assign addr[3742]= 2090184478;
assign addr[3743]= 2106406677;
assign addr[3744]= 2119956737;
assign addr[3745]= 2130817471;
assign addr[3746]= 2138975100;
assign addr[3747]= 2144419275;
assign addr[3748]= 2147143090;
assign addr[3749]= 2147143090;
assign addr[3750]= 2144419275;
assign addr[3751]= 2138975100;
assign addr[3752]= 2130817471;
assign addr[3753]= 2119956737;
assign addr[3754]= 2106406677;
assign addr[3755]= 2090184478;
assign addr[3756]= 2071310720;
assign addr[3757]= 2049809346;
assign addr[3758]= 2025707632;
assign addr[3759]= 1999036154;
assign addr[3760]= 1969828744;
assign addr[3761]= 1938122457;
assign addr[3762]= 1903957513;
assign addr[3763]= 1867377253;
assign addr[3764]= 1828428082;
assign addr[3765]= 1787159411;
assign addr[3766]= 1743623590;
assign addr[3767]= 1697875851;
assign addr[3768]= 1649974225;
assign addr[3769]= 1599979481;
assign addr[3770]= 1547955041;
assign addr[3771]= 1493966902;
assign addr[3772]= 1438083551;
assign addr[3773]= 1380375881;
assign addr[3774]= 1320917099;
assign addr[3775]= 1259782632;
assign addr[3776]= 1197050035;
assign addr[3777]= 1132798888;
assign addr[3778]= 1067110699;
assign addr[3779]= 1000068799;
assign addr[3780]= 931758235;
assign addr[3781]= 862265664;
assign addr[3782]= 791679244;
assign addr[3783]= 720088517;
assign addr[3784]= 647584304;
assign addr[3785]= 574258580;
assign addr[3786]= 500204365;
assign addr[3787]= 425515602;
assign addr[3788]= 350287041;
assign addr[3789]= 274614114;
assign addr[3790]= 198592817;
assign addr[3791]= 122319591;
assign addr[3792]= 45891193;
assign addr[3793]= -30595422;
assign addr[3794]= -107043224;
assign addr[3795]= -183355234;
assign addr[3796]= -259434643;
assign addr[3797]= -335184940;
assign addr[3798]= -410510029;
assign addr[3799]= -485314355;
assign addr[3800]= -559503022;
assign addr[3801]= -632981917;
assign addr[3802]= -705657826;
assign addr[3803]= -777438554;
assign addr[3804]= -848233042;
assign addr[3805]= -917951481;
assign addr[3806]= -986505429;
assign addr[3807]= -1053807919;
assign addr[3808]= -1119773573;
assign addr[3809]= -1184318708;
assign addr[3810]= -1247361445;
assign addr[3811]= -1308821808;
assign addr[3812]= -1368621831;
assign addr[3813]= -1426685652;
assign addr[3814]= -1482939614;
assign addr[3815]= -1537312353;
assign addr[3816]= -1589734894;
assign addr[3817]= -1640140734;
assign addr[3818]= -1688465931;
assign addr[3819]= -1734649179;
assign addr[3820]= -1778631892;
assign addr[3821]= -1820358275;
assign addr[3822]= -1859775393;
assign addr[3823]= -1896833245;
assign addr[3824]= -1931484818;
assign addr[3825]= -1963686155;
assign addr[3826]= -1993396407;
assign addr[3827]= -2020577882;
assign addr[3828]= -2045196100;
assign addr[3829]= -2067219829;
assign addr[3830]= -2086621133;
assign addr[3831]= -2103375398;
assign addr[3832]= -2117461370;
assign addr[3833]= -2128861181;
assign addr[3834]= -2137560369;
assign addr[3835]= -2143547897;
assign addr[3836]= -2146816171;
assign addr[3837]= -2147361045;
assign addr[3838]= -2145181827;
assign addr[3839]= -2140281282;
assign addr[3840]= -2132665626;
assign addr[3841]= -2122344521;
assign addr[3842]= -2109331059;
assign addr[3843]= -2093641749;
assign addr[3844]= -2075296495;
assign addr[3845]= -2054318569;
assign addr[3846]= -2030734582;
assign addr[3847]= -2004574453;
assign addr[3848]= -1975871368;
assign addr[3849]= -1944661739;
assign addr[3850]= -1910985158;
assign addr[3851]= -1874884346;
assign addr[3852]= -1836405100;
assign addr[3853]= -1795596234;
assign addr[3854]= -1752509516;
assign addr[3855]= -1707199606;
assign addr[3856]= -1659723983;
assign addr[3857]= -1610142873;
assign addr[3858]= -1558519173;
assign addr[3859]= -1504918373;
assign addr[3860]= -1449408469;
assign addr[3861]= -1392059879;
assign addr[3862]= -1332945355;
assign addr[3863]= -1272139887;
assign addr[3864]= -1209720613;
assign addr[3865]= -1145766716;
assign addr[3866]= -1080359326;
assign addr[3867]= -1013581418;
assign addr[3868]= -945517704;
assign addr[3869]= -876254528;
assign addr[3870]= -805879757;
assign addr[3871]= -734482665;
assign addr[3872]= -662153826;
assign addr[3873]= -588984994;
assign addr[3874]= -515068990;
assign addr[3875]= -440499581;
assign addr[3876]= -365371365;
assign addr[3877]= -289779648;
assign addr[3878]= -213820322;
assign addr[3879]= -137589750;
assign addr[3880]= -61184634;
assign addr[3881]= 15298099;
assign addr[3882]= 91761426;
assign addr[3883]= 168108346;
assign addr[3884]= 244242007;
assign addr[3885]= 320065829;
assign addr[3886]= 395483624;
assign addr[3887]= 470399716;
assign addr[3888]= 544719071;
assign addr[3889]= 618347408;
assign addr[3890]= 691191324;
assign addr[3891]= 763158411;
assign addr[3892]= 834157373;
assign addr[3893]= 904098143;
assign addr[3894]= 972891995;
assign addr[3895]= 1040451659;
assign addr[3896]= 1106691431;
assign addr[3897]= 1171527280;
assign addr[3898]= 1234876957;
assign addr[3899]= 1296660098;
assign addr[3900]= 1356798326;
assign addr[3901]= 1415215352;
assign addr[3902]= 1471837070;
assign addr[3903]= 1526591649;
assign addr[3904]= 1579409630;
assign addr[3905]= 1630224009;
assign addr[3906]= 1678970324;
assign addr[3907]= 1725586737;
assign addr[3908]= 1770014111;
assign addr[3909]= 1812196087;
assign addr[3910]= 1852079154;
assign addr[3911]= 1889612716;
assign addr[3912]= 1924749160;
assign addr[3913]= 1957443913;
assign addr[3914]= 1987655498;
assign addr[3915]= 2015345591;
assign addr[3916]= 2040479063;
assign addr[3917]= 2063024031;
assign addr[3918]= 2082951896;
assign addr[3919]= 2100237377;
assign addr[3920]= 2114858546;
assign addr[3921]= 2126796855;
assign addr[3922]= 2136037160;
assign addr[3923]= 2142567738;
assign addr[3924]= 2146380306;
assign addr[3925]= 2147470025;
assign addr[3926]= 2145835515;
assign addr[3927]= 2141478848;
assign addr[3928]= 2134405552;
assign addr[3929]= 2124624598;
assign addr[3930]= 2112148396;
assign addr[3931]= 2096992772;
assign addr[3932]= 2079176953;
assign addr[3933]= 2058723538;
assign addr[3934]= 2035658475;
assign addr[3935]= 2010011024;
assign addr[3936]= 1981813720;
assign addr[3937]= 1951102334;
assign addr[3938]= 1917915825;
assign addr[3939]= 1882296293;
assign addr[3940]= 1844288924;
assign addr[3941]= 1803941934;
assign addr[3942]= 1761306505;
assign addr[3943]= 1716436725;
assign addr[3944]= 1669389513;
assign addr[3945]= 1620224553;
assign addr[3946]= 1569004214;
assign addr[3947]= 1515793473;
assign addr[3948]= 1460659832;
assign addr[3949]= 1403673233;
assign addr[3950]= 1344905966;
assign addr[3951]= 1284432584;
assign addr[3952]= 1222329801;
assign addr[3953]= 1158676398;
assign addr[3954]= 1093553126;
assign addr[3955]= 1027042599;
assign addr[3956]= 959229189;
assign addr[3957]= 890198924;
assign addr[3958]= 820039373;
assign addr[3959]= 748839539;
assign addr[3960]= 676689746;
assign addr[3961]= 603681519;
assign addr[3962]= 529907477;
assign addr[3963]= 455461206;
assign addr[3964]= 380437148;
assign addr[3965]= 304930476;
assign addr[3966]= 229036977;
assign addr[3967]= 152852926;
assign addr[3968]= 76474970;
assign addr[3969]= 0;
assign addr[3970]= -76474970;
assign addr[3971]= -152852926;
assign addr[3972]= -229036977;
assign addr[3973]= -304930476;
assign addr[3974]= -380437148;
assign addr[3975]= -455461206;
assign addr[3976]= -529907477;
assign addr[3977]= -603681519;
assign addr[3978]= -676689746;
assign addr[3979]= -748839539;
assign addr[3980]= -820039373;
assign addr[3981]= -890198924;
assign addr[3982]= -959229189;
assign addr[3983]= -1027042599;
assign addr[3984]= -1093553126;
assign addr[3985]= -1158676398;
assign addr[3986]= -1222329801;
assign addr[3987]= -1284432584;
assign addr[3988]= -1344905966;
assign addr[3989]= -1403673233;
assign addr[3990]= -1460659832;
assign addr[3991]= -1515793473;
assign addr[3992]= -1569004214;
assign addr[3993]= -1620224553;
assign addr[3994]= -1669389513;
assign addr[3995]= -1716436725;
assign addr[3996]= -1761306505;
assign addr[3997]= -1803941934;
assign addr[3998]= -1844288924;
assign addr[3999]= -1882296293;
assign addr[4000]= -1917915825;
assign addr[4001]= -1951102334;
assign addr[4002]= -1981813720;
assign addr[4003]= -2010011024;
assign addr[4004]= -2035658475;
assign addr[4005]= -2058723538;
assign addr[4006]= -2079176953;
assign addr[4007]= -2096992772;
assign addr[4008]= -2112148396;
assign addr[4009]= -2124624598;
assign addr[4010]= -2134405552;
assign addr[4011]= -2141478848;
assign addr[4012]= -2145835515;
assign addr[4013]= -2147470025;
assign addr[4014]= -2146380306;
assign addr[4015]= -2142567738;
assign addr[4016]= -2136037160;
assign addr[4017]= -2126796855;
assign addr[4018]= -2114858546;
assign addr[4019]= -2100237377;
assign addr[4020]= -2082951896;
assign addr[4021]= -2063024031;
assign addr[4022]= -2040479063;
assign addr[4023]= -2015345591;
assign addr[4024]= -1987655498;
assign addr[4025]= -1957443913;
assign addr[4026]= -1924749160;
assign addr[4027]= -1889612716;
assign addr[4028]= -1852079154;
assign addr[4029]= -1812196087;
assign addr[4030]= -1770014111;
assign addr[4031]= -1725586737;
assign addr[4032]= -1678970324;
assign addr[4033]= -1630224009;
assign addr[4034]= -1579409630;
assign addr[4035]= -1526591649;
assign addr[4036]= -1471837070;
assign addr[4037]= -1415215352;
assign addr[4038]= -1356798326;
assign addr[4039]= -1296660098;
assign addr[4040]= -1234876957;
assign addr[4041]= -1171527280;
assign addr[4042]= -1106691431;
assign addr[4043]= -1040451659;
assign addr[4044]= -972891995;
assign addr[4045]= -904098143;
assign addr[4046]= -834157373;
assign addr[4047]= -763158411;
assign addr[4048]= -691191324;
assign addr[4049]= -618347408;
assign addr[4050]= -544719071;
assign addr[4051]= -470399716;
assign addr[4052]= -395483624;
assign addr[4053]= -320065829;
assign addr[4054]= -244242007;
assign addr[4055]= -168108346;
assign addr[4056]= -91761426;
assign addr[4057]= -15298099;
assign addr[4058]= 61184634;
assign addr[4059]= 137589750;
assign addr[4060]= 213820322;
assign addr[4061]= 289779648;
assign addr[4062]= 365371365;
assign addr[4063]= 440499581;
assign addr[4064]= 515068990;
assign addr[4065]= 588984994;
assign addr[4066]= 662153826;
assign addr[4067]= 734482665;
assign addr[4068]= 805879757;
assign addr[4069]= 876254528;
assign addr[4070]= 945517704;
assign addr[4071]= 1013581418;
assign addr[4072]= 1080359326;
assign addr[4073]= 1145766716;
assign addr[4074]= 1209720613;
assign addr[4075]= 1272139887;
assign addr[4076]= 1332945355;
assign addr[4077]= 1392059879;
assign addr[4078]= 1449408469;
assign addr[4079]= 1504918373;
assign addr[4080]= 1558519173;
assign addr[4081]= 1610142873;
assign addr[4082]= 1659723983;
assign addr[4083]= 1707199606;
assign addr[4084]= 1752509516;
assign addr[4085]= 1795596234;
assign addr[4086]= 1836405100;
assign addr[4087]= 1874884346;
assign addr[4088]= 1910985158;
assign addr[4089]= 1944661739;
assign addr[4090]= 1975871368;
assign addr[4091]= 2004574453;
assign addr[4092]= 2030734582;
assign addr[4093]= 2054318569;
assign addr[4094]= 2075296495;
assign addr[4095]= 2093641749;
assign addr[4096]= 2109331059;
assign addr[4097]= 2122344521;
assign addr[4098]= 2132665626;
assign addr[4099]= 2140281282;
assign addr[4100]= 2145181827;
assign addr[4101]= 2147361045;
assign addr[4102]= 2146816171;
assign addr[4103]= 2143547897;
assign addr[4104]= 2137560369;
assign addr[4105]= 2128861181;
assign addr[4106]= 2117461370;
assign addr[4107]= 2103375398;
assign addr[4108]= 2086621133;
assign addr[4109]= 2067219829;
assign addr[4110]= 2045196100;
assign addr[4111]= 2020577882;
assign addr[4112]= 1993396407;
assign addr[4113]= 1963686155;
assign addr[4114]= 1931484818;
assign addr[4115]= 1896833245;
assign addr[4116]= 1859775393;
assign addr[4117]= 1820358275;
assign addr[4118]= 1778631892;
assign addr[4119]= 1734649179;
assign addr[4120]= 1688465931;
assign addr[4121]= 1640140734;
assign addr[4122]= 1589734894;
assign addr[4123]= 1537312353;
assign addr[4124]= 1482939614;
assign addr[4125]= 1426685652;
assign addr[4126]= 1368621831;
assign addr[4127]= 1308821808;
assign addr[4128]= 1247361445;
assign addr[4129]= 1184318708;
assign addr[4130]= 1119773573;
assign addr[4131]= 1053807919;
assign addr[4132]= 986505429;
assign addr[4133]= 917951481;
assign addr[4134]= 848233042;
assign addr[4135]= 777438554;
assign addr[4136]= 705657826;
assign addr[4137]= 632981917;
assign addr[4138]= 559503022;
assign addr[4139]= 485314355;
assign addr[4140]= 410510029;
assign addr[4141]= 335184940;
assign addr[4142]= 259434643;
assign addr[4143]= 183355234;
assign addr[4144]= 107043224;
assign addr[4145]= 30595422;
assign addr[4146]= -45891193;
assign addr[4147]= -122319591;
assign addr[4148]= -198592817;
assign addr[4149]= -274614114;
assign addr[4150]= -350287041;
assign addr[4151]= -425515602;
assign addr[4152]= -500204365;
assign addr[4153]= -574258580;
assign addr[4154]= -647584304;
assign addr[4155]= -720088517;
assign addr[4156]= -791679244;
assign addr[4157]= -862265664;
assign addr[4158]= -931758235;
assign addr[4159]= -1000068799;
assign addr[4160]= -1067110699;
assign addr[4161]= -1132798888;
assign addr[4162]= -1197050035;
assign addr[4163]= -1259782632;
assign addr[4164]= -1320917099;
assign addr[4165]= -1380375881;
assign addr[4166]= -1438083551;
assign addr[4167]= -1493966902;
assign addr[4168]= -1547955041;
assign addr[4169]= -1599979481;
assign addr[4170]= -1649974225;
assign addr[4171]= -1697875851;
assign addr[4172]= -1743623590;
assign addr[4173]= -1787159411;
assign addr[4174]= -1828428082;
assign addr[4175]= -1867377253;
assign addr[4176]= -1903957513;
assign addr[4177]= -1938122457;
assign addr[4178]= -1969828744;
assign addr[4179]= -1999036154;
assign addr[4180]= -2025707632;
assign addr[4181]= -2049809346;
assign addr[4182]= -2071310720;
assign addr[4183]= -2090184478;
assign addr[4184]= -2106406677;
assign addr[4185]= -2119956737;
assign addr[4186]= -2130817471;
assign addr[4187]= -2138975100;
assign addr[4188]= -2144419275;
assign addr[4189]= -2147143090;
assign addr[4190]= -2147143090;
assign addr[4191]= -2144419275;
assign addr[4192]= -2138975100;
assign addr[4193]= -2130817471;
assign addr[4194]= -2119956737;
assign addr[4195]= -2106406677;
assign addr[4196]= -2090184478;
assign addr[4197]= -2071310720;
assign addr[4198]= -2049809346;
assign addr[4199]= -2025707632;
assign addr[4200]= -1999036154;
assign addr[4201]= -1969828744;
assign addr[4202]= -1938122457;
assign addr[4203]= -1903957513;
assign addr[4204]= -1867377253;
assign addr[4205]= -1828428082;
assign addr[4206]= -1787159411;
assign addr[4207]= -1743623590;
assign addr[4208]= -1697875851;
assign addr[4209]= -1649974225;
assign addr[4210]= -1599979481;
assign addr[4211]= -1547955041;
assign addr[4212]= -1493966902;
assign addr[4213]= -1438083551;
assign addr[4214]= -1380375881;
assign addr[4215]= -1320917099;
assign addr[4216]= -1259782632;
assign addr[4217]= -1197050035;
assign addr[4218]= -1132798888;
assign addr[4219]= -1067110699;
assign addr[4220]= -1000068799;
assign addr[4221]= -931758235;
assign addr[4222]= -862265664;
assign addr[4223]= -791679244;
assign addr[4224]= -720088517;
assign addr[4225]= -647584304;
assign addr[4226]= -574258580;
assign addr[4227]= -500204365;
assign addr[4228]= -425515602;
assign addr[4229]= -350287041;
assign addr[4230]= -274614114;
assign addr[4231]= -198592817;
assign addr[4232]= -122319591;
assign addr[4233]= -45891193;
assign addr[4234]= 30595422;
assign addr[4235]= 107043224;
assign addr[4236]= 183355234;
assign addr[4237]= 259434643;
assign addr[4238]= 335184940;
assign addr[4239]= 410510029;
assign addr[4240]= 485314355;
assign addr[4241]= 559503022;
assign addr[4242]= 632981917;
assign addr[4243]= 705657826;
assign addr[4244]= 777438554;
assign addr[4245]= 848233042;
assign addr[4246]= 917951481;
assign addr[4247]= 986505429;
assign addr[4248]= 1053807919;
assign addr[4249]= 1119773573;
assign addr[4250]= 1184318708;
assign addr[4251]= 1247361445;
assign addr[4252]= 1308821808;
assign addr[4253]= 1368621831;
assign addr[4254]= 1426685652;
assign addr[4255]= 1482939614;
assign addr[4256]= 1537312353;
assign addr[4257]= 1589734894;
assign addr[4258]= 1640140734;
assign addr[4259]= 1688465931;
assign addr[4260]= 1734649179;
assign addr[4261]= 1778631892;
assign addr[4262]= 1820358275;
assign addr[4263]= 1859775393;
assign addr[4264]= 1896833245;
assign addr[4265]= 1931484818;
assign addr[4266]= 1963686155;
assign addr[4267]= 1993396407;
assign addr[4268]= 2020577882;
assign addr[4269]= 2045196100;
assign addr[4270]= 2067219829;
assign addr[4271]= 2086621133;
assign addr[4272]= 2103375398;
assign addr[4273]= 2117461370;
assign addr[4274]= 2128861181;
assign addr[4275]= 2137560369;
assign addr[4276]= 2143547897;
assign addr[4277]= 2146816171;
assign addr[4278]= 2147361045;
assign addr[4279]= 2145181827;
assign addr[4280]= 2140281282;
assign addr[4281]= 2132665626;
assign addr[4282]= 2122344521;
assign addr[4283]= 2109331059;
assign addr[4284]= 2093641749;
assign addr[4285]= 2075296495;
assign addr[4286]= 2054318569;
assign addr[4287]= 2030734582;
assign addr[4288]= 2004574453;
assign addr[4289]= 1975871368;
assign addr[4290]= 1944661739;
assign addr[4291]= 1910985158;
assign addr[4292]= 1874884346;
assign addr[4293]= 1836405100;
assign addr[4294]= 1795596234;
assign addr[4295]= 1752509516;
assign addr[4296]= 1707199606;
assign addr[4297]= 1659723983;
assign addr[4298]= 1610142873;
assign addr[4299]= 1558519173;
assign addr[4300]= 1504918373;
assign addr[4301]= 1449408469;
assign addr[4302]= 1392059879;
assign addr[4303]= 1332945355;
assign addr[4304]= 1272139887;
assign addr[4305]= 1209720613;
assign addr[4306]= 1145766716;
assign addr[4307]= 1080359326;
assign addr[4308]= 1013581418;
assign addr[4309]= 945517704;
assign addr[4310]= 876254528;
assign addr[4311]= 805879757;
assign addr[4312]= 734482665;
assign addr[4313]= 662153826;
assign addr[4314]= 588984994;
assign addr[4315]= 515068990;
assign addr[4316]= 440499581;
assign addr[4317]= 365371365;
assign addr[4318]= 289779648;
assign addr[4319]= 213820322;
assign addr[4320]= 137589750;
assign addr[4321]= 61184634;
assign addr[4322]= -15298099;
assign addr[4323]= -91761426;
assign addr[4324]= -168108346;
assign addr[4325]= -244242007;
assign addr[4326]= -320065829;
assign addr[4327]= -395483624;
assign addr[4328]= -470399716;
assign addr[4329]= -544719071;
assign addr[4330]= -618347408;
assign addr[4331]= -691191324;
assign addr[4332]= -763158411;
assign addr[4333]= -834157373;
assign addr[4334]= -904098143;
assign addr[4335]= -972891995;
assign addr[4336]= -1040451659;
assign addr[4337]= -1106691431;
assign addr[4338]= -1171527280;
assign addr[4339]= -1234876957;
assign addr[4340]= -1296660098;
assign addr[4341]= -1356798326;
assign addr[4342]= -1415215352;
assign addr[4343]= -1471837070;
assign addr[4344]= -1526591649;
assign addr[4345]= -1579409630;
assign addr[4346]= -1630224009;
assign addr[4347]= -1678970324;
assign addr[4348]= -1725586737;
assign addr[4349]= -1770014111;
assign addr[4350]= -1812196087;
assign addr[4351]= -1852079154;
assign addr[4352]= -1889612716;
assign addr[4353]= -1924749160;
assign addr[4354]= -1957443913;
assign addr[4355]= -1987655498;
assign addr[4356]= -2015345591;
assign addr[4357]= -2040479063;
assign addr[4358]= -2063024031;
assign addr[4359]= -2082951896;
assign addr[4360]= -2100237377;
assign addr[4361]= -2114858546;
assign addr[4362]= -2126796855;
assign addr[4363]= -2136037160;
assign addr[4364]= -2142567738;
assign addr[4365]= -2146380306;
assign addr[4366]= -2147470025;
assign addr[4367]= -2145835515;
assign addr[4368]= -2141478848;
assign addr[4369]= -2134405552;
assign addr[4370]= -2124624598;
assign addr[4371]= -2112148396;
assign addr[4372]= -2096992772;
assign addr[4373]= -2079176953;
assign addr[4374]= -2058723538;
assign addr[4375]= -2035658475;
assign addr[4376]= -2010011024;
assign addr[4377]= -1981813720;
assign addr[4378]= -1951102334;
assign addr[4379]= -1917915825;
assign addr[4380]= -1882296293;
assign addr[4381]= -1844288924;
assign addr[4382]= -1803941934;
assign addr[4383]= -1761306505;
assign addr[4384]= -1716436725;
assign addr[4385]= -1669389513;
assign addr[4386]= -1620224553;
assign addr[4387]= -1569004214;
assign addr[4388]= -1515793473;
assign addr[4389]= -1460659832;
assign addr[4390]= -1403673233;
assign addr[4391]= -1344905966;
assign addr[4392]= -1284432584;
assign addr[4393]= -1222329801;
assign addr[4394]= -1158676398;
assign addr[4395]= -1093553126;
assign addr[4396]= -1027042599;
assign addr[4397]= -959229189;
assign addr[4398]= -890198924;
assign addr[4399]= -820039373;
assign addr[4400]= -748839539;
assign addr[4401]= -676689746;
assign addr[4402]= -603681519;
assign addr[4403]= -529907477;
assign addr[4404]= -455461206;
assign addr[4405]= -380437148;
assign addr[4406]= -304930476;
assign addr[4407]= -229036977;
assign addr[4408]= -152852926;
assign addr[4409]= -76474970;
assign addr[4410]= 0;
assign addr[4411]= 76474970;
assign addr[4412]= 152852926;
assign addr[4413]= 229036977;
assign addr[4414]= 304930476;
assign addr[4415]= 380437148;
assign addr[4416]= 455461206;
assign addr[4417]= 529907477;
assign addr[4418]= 603681519;
assign addr[4419]= 676689746;
assign addr[4420]= 748839539;
assign addr[4421]= 820039373;
assign addr[4422]= 890198924;
assign addr[4423]= 959229189;
assign addr[4424]= 1027042599;
assign addr[4425]= 1093553126;
assign addr[4426]= 1158676398;
assign addr[4427]= 1222329801;
assign addr[4428]= 1284432584;
assign addr[4429]= 1344905966;
assign addr[4430]= 1403673233;
assign addr[4431]= 1460659832;
assign addr[4432]= 1515793473;
assign addr[4433]= 1569004214;
assign addr[4434]= 1620224553;
assign addr[4435]= 1669389513;
assign addr[4436]= 1716436725;
assign addr[4437]= 1761306505;
assign addr[4438]= 1803941934;
assign addr[4439]= 1844288924;
assign addr[4440]= 1882296293;
assign addr[4441]= 1917915825;
assign addr[4442]= 1951102334;
assign addr[4443]= 1981813720;
assign addr[4444]= 2010011024;
assign addr[4445]= 2035658475;
assign addr[4446]= 2058723538;
assign addr[4447]= 2079176953;
assign addr[4448]= 2096992772;
assign addr[4449]= 2112148396;
assign addr[4450]= 2124624598;
assign addr[4451]= 2134405552;
assign addr[4452]= 2141478848;
assign addr[4453]= 2145835515;
assign addr[4454]= 2147470025;
assign addr[4455]= 2146380306;
assign addr[4456]= 2142567738;
assign addr[4457]= 2136037160;
assign addr[4458]= 2126796855;
assign addr[4459]= 2114858546;
assign addr[4460]= 2100237377;
assign addr[4461]= 2082951896;
assign addr[4462]= 2063024031;
assign addr[4463]= 2040479063;
assign addr[4464]= 2015345591;
assign addr[4465]= 1987655498;
assign addr[4466]= 1957443913;
assign addr[4467]= 1924749160;
assign addr[4468]= 1889612716;
assign addr[4469]= 1852079154;
assign addr[4470]= 1812196087;
assign addr[4471]= 1770014111;
assign addr[4472]= 1725586737;
assign addr[4473]= 1678970324;
assign addr[4474]= 1630224009;
assign addr[4475]= 1579409630;
assign addr[4476]= 1526591649;
assign addr[4477]= 1471837070;
assign addr[4478]= 1415215352;
assign addr[4479]= 1356798326;
assign addr[4480]= 1296660098;
assign addr[4481]= 1234876957;
assign addr[4482]= 1171527280;
assign addr[4483]= 1106691431;
assign addr[4484]= 1040451659;
assign addr[4485]= 972891995;
assign addr[4486]= 904098143;
assign addr[4487]= 834157373;
assign addr[4488]= 763158411;
assign addr[4489]= 691191324;
assign addr[4490]= 618347408;
assign addr[4491]= 544719071;
assign addr[4492]= 470399716;
assign addr[4493]= 395483624;
assign addr[4494]= 320065829;
assign addr[4495]= 244242007;
assign addr[4496]= 168108346;
assign addr[4497]= 91761426;
assign addr[4498]= 15298099;
assign addr[4499]= -61184634;
assign addr[4500]= -137589750;
assign addr[4501]= -213820322;
assign addr[4502]= -289779648;
assign addr[4503]= -365371365;
assign addr[4504]= -440499581;
assign addr[4505]= -515068990;
assign addr[4506]= -588984994;
assign addr[4507]= -662153826;
assign addr[4508]= -734482665;
assign addr[4509]= -805879757;
assign addr[4510]= -876254528;
assign addr[4511]= -945517704;
assign addr[4512]= -1013581418;
assign addr[4513]= -1080359326;
assign addr[4514]= -1145766716;
assign addr[4515]= -1209720613;
assign addr[4516]= -1272139887;
assign addr[4517]= -1332945355;
assign addr[4518]= -1392059879;
assign addr[4519]= -1449408469;
assign addr[4520]= -1504918373;
assign addr[4521]= -1558519173;
assign addr[4522]= -1610142873;
assign addr[4523]= -1659723983;
assign addr[4524]= -1707199606;
assign addr[4525]= -1752509516;
assign addr[4526]= -1795596234;
assign addr[4527]= -1836405100;
assign addr[4528]= -1874884346;
assign addr[4529]= -1910985158;
assign addr[4530]= -1944661739;
assign addr[4531]= -1975871368;
assign addr[4532]= -2004574453;
assign addr[4533]= -2030734582;
assign addr[4534]= -2054318569;
assign addr[4535]= -2075296495;
assign addr[4536]= -2093641749;
assign addr[4537]= -2109331059;
assign addr[4538]= -2122344521;
assign addr[4539]= -2132665626;
assign addr[4540]= -2140281282;
assign addr[4541]= -2145181827;
assign addr[4542]= -2147361045;
assign addr[4543]= -2146816171;
assign addr[4544]= -2143547897;
assign addr[4545]= -2137560369;
assign addr[4546]= -2128861181;
assign addr[4547]= -2117461370;
assign addr[4548]= -2103375398;
assign addr[4549]= -2086621133;
assign addr[4550]= -2067219829;
assign addr[4551]= -2045196100;
assign addr[4552]= -2020577882;
assign addr[4553]= -1993396407;
assign addr[4554]= -1963686155;
assign addr[4555]= -1931484818;
assign addr[4556]= -1896833245;
assign addr[4557]= -1859775393;
assign addr[4558]= -1820358275;
assign addr[4559]= -1778631892;
assign addr[4560]= -1734649179;
assign addr[4561]= -1688465931;
assign addr[4562]= -1640140734;
assign addr[4563]= -1589734894;
assign addr[4564]= -1537312353;
assign addr[4565]= -1482939614;
assign addr[4566]= -1426685652;
assign addr[4567]= -1368621831;
assign addr[4568]= -1308821808;
assign addr[4569]= -1247361445;
assign addr[4570]= -1184318708;
assign addr[4571]= -1119773573;
assign addr[4572]= -1053807919;
assign addr[4573]= -986505429;
assign addr[4574]= -917951481;
assign addr[4575]= -848233042;
assign addr[4576]= -777438554;
assign addr[4577]= -705657826;
assign addr[4578]= -632981917;
assign addr[4579]= -559503022;
assign addr[4580]= -485314355;
assign addr[4581]= -410510029;
assign addr[4582]= -335184940;
assign addr[4583]= -259434643;
assign addr[4584]= -183355234;
assign addr[4585]= -107043224;
assign addr[4586]= -30595422;
assign addr[4587]= 45891193;
assign addr[4588]= 122319591;
assign addr[4589]= 198592817;
assign addr[4590]= 274614114;
assign addr[4591]= 350287041;
assign addr[4592]= 425515602;
assign addr[4593]= 500204365;
assign addr[4594]= 574258580;
assign addr[4595]= 647584304;
assign addr[4596]= 720088517;
assign addr[4597]= 791679244;
assign addr[4598]= 862265664;
assign addr[4599]= 931758235;
assign addr[4600]= 1000068799;
assign addr[4601]= 1067110699;
assign addr[4602]= 1132798888;
assign addr[4603]= 1197050035;
assign addr[4604]= 1259782632;
assign addr[4605]= 1320917099;
assign addr[4606]= 1380375881;
assign addr[4607]= 1438083551;
assign addr[4608]= 1493966902;
assign addr[4609]= 1547955041;
assign addr[4610]= 1599979481;
assign addr[4611]= 1649974225;
assign addr[4612]= 1697875851;
assign addr[4613]= 1743623590;
assign addr[4614]= 1787159411;
assign addr[4615]= 1828428082;
assign addr[4616]= 1867377253;
assign addr[4617]= 1903957513;
assign addr[4618]= 1938122457;
assign addr[4619]= 1969828744;
assign addr[4620]= 1999036154;
assign addr[4621]= 2025707632;
assign addr[4622]= 2049809346;
assign addr[4623]= 2071310720;
assign addr[4624]= 2090184478;
assign addr[4625]= 2106406677;
assign addr[4626]= 2119956737;
assign addr[4627]= 2130817471;
assign addr[4628]= 2138975100;
assign addr[4629]= 2144419275;
assign addr[4630]= 2147143090;
assign addr[4631]= 2147143090;
assign addr[4632]= 2144419275;
assign addr[4633]= 2138975100;
assign addr[4634]= 2130817471;
assign addr[4635]= 2119956737;
assign addr[4636]= 2106406677;
assign addr[4637]= 2090184478;
assign addr[4638]= 2071310720;
assign addr[4639]= 2049809346;
assign addr[4640]= 2025707632;
assign addr[4641]= 1999036154;
assign addr[4642]= 1969828744;
assign addr[4643]= 1938122457;
assign addr[4644]= 1903957513;
assign addr[4645]= 1867377253;
assign addr[4646]= 1828428082;
assign addr[4647]= 1787159411;
assign addr[4648]= 1743623590;
assign addr[4649]= 1697875851;
assign addr[4650]= 1649974225;
assign addr[4651]= 1599979481;
assign addr[4652]= 1547955041;
assign addr[4653]= 1493966902;
assign addr[4654]= 1438083551;
assign addr[4655]= 1380375881;
assign addr[4656]= 1320917099;
assign addr[4657]= 1259782632;
assign addr[4658]= 1197050035;
assign addr[4659]= 1132798888;
assign addr[4660]= 1067110699;
assign addr[4661]= 1000068799;
assign addr[4662]= 931758235;
assign addr[4663]= 862265664;
assign addr[4664]= 791679244;
assign addr[4665]= 720088517;
assign addr[4666]= 647584304;
assign addr[4667]= 574258580;
assign addr[4668]= 500204365;
assign addr[4669]= 425515602;
assign addr[4670]= 350287041;
assign addr[4671]= 274614114;
assign addr[4672]= 198592817;
assign addr[4673]= 122319591;
assign addr[4674]= 45891193;
assign addr[4675]= -30595422;
assign addr[4676]= -107043224;
assign addr[4677]= -183355234;
assign addr[4678]= -259434643;
assign addr[4679]= -335184940;
assign addr[4680]= -410510029;
assign addr[4681]= -485314355;
assign addr[4682]= -559503022;
assign addr[4683]= -632981917;
assign addr[4684]= -705657826;
assign addr[4685]= -777438554;
assign addr[4686]= -848233042;
assign addr[4687]= -917951481;
assign addr[4688]= -986505429;
assign addr[4689]= -1053807919;
assign addr[4690]= -1119773573;
assign addr[4691]= -1184318708;
assign addr[4692]= -1247361445;
assign addr[4693]= -1308821808;
assign addr[4694]= -1368621831;
assign addr[4695]= -1426685652;
assign addr[4696]= -1482939614;
assign addr[4697]= -1537312353;
assign addr[4698]= -1589734894;
assign addr[4699]= -1640140734;
assign addr[4700]= -1688465931;
assign addr[4701]= -1734649179;
assign addr[4702]= -1778631892;
assign addr[4703]= -1820358275;
assign addr[4704]= -1859775393;
assign addr[4705]= -1896833245;
assign addr[4706]= -1931484818;
assign addr[4707]= -1963686155;
assign addr[4708]= -1993396407;
assign addr[4709]= -2020577882;
assign addr[4710]= -2045196100;
assign addr[4711]= -2067219829;
assign addr[4712]= -2086621133;
assign addr[4713]= -2103375398;
assign addr[4714]= -2117461370;
assign addr[4715]= -2128861181;
assign addr[4716]= -2137560369;
assign addr[4717]= -2143547897;
assign addr[4718]= -2146816171;
assign addr[4719]= -2147361045;
assign addr[4720]= -2145181827;
assign addr[4721]= -2140281282;
assign addr[4722]= -2132665626;
assign addr[4723]= -2122344521;
assign addr[4724]= -2109331059;
assign addr[4725]= -2093641749;
assign addr[4726]= -2075296495;
assign addr[4727]= -2054318569;
assign addr[4728]= -2030734582;
assign addr[4729]= -2004574453;
assign addr[4730]= -1975871368;
assign addr[4731]= -1944661739;
assign addr[4732]= -1910985158;
assign addr[4733]= -1874884346;
assign addr[4734]= -1836405100;
assign addr[4735]= -1795596234;
assign addr[4736]= -1752509516;
assign addr[4737]= -1707199606;
assign addr[4738]= -1659723983;
assign addr[4739]= -1610142873;
assign addr[4740]= -1558519173;
assign addr[4741]= -1504918373;
assign addr[4742]= -1449408469;
assign addr[4743]= -1392059879;
assign addr[4744]= -1332945355;
assign addr[4745]= -1272139887;
assign addr[4746]= -1209720613;
assign addr[4747]= -1145766716;
assign addr[4748]= -1080359326;
assign addr[4749]= -1013581418;
assign addr[4750]= -945517704;
assign addr[4751]= -876254528;
assign addr[4752]= -805879757;
assign addr[4753]= -734482665;
assign addr[4754]= -662153826;
assign addr[4755]= -588984994;
assign addr[4756]= -515068990;
assign addr[4757]= -440499581;
assign addr[4758]= -365371365;
assign addr[4759]= -289779648;
assign addr[4760]= -213820322;
assign addr[4761]= -137589750;
assign addr[4762]= -61184634;
assign addr[4763]= 15298099;
assign addr[4764]= 91761426;
assign addr[4765]= 168108346;
assign addr[4766]= 244242007;
assign addr[4767]= 320065829;
assign addr[4768]= 395483624;
assign addr[4769]= 470399716;
assign addr[4770]= 544719071;
assign addr[4771]= 618347408;
assign addr[4772]= 691191324;
assign addr[4773]= 763158411;
assign addr[4774]= 834157373;
assign addr[4775]= 904098143;
assign addr[4776]= 972891995;
assign addr[4777]= 1040451659;
assign addr[4778]= 1106691431;
assign addr[4779]= 1171527280;
assign addr[4780]= 1234876957;
assign addr[4781]= 1296660098;
assign addr[4782]= 1356798326;
assign addr[4783]= 1415215352;
assign addr[4784]= 1471837070;
assign addr[4785]= 1526591649;
assign addr[4786]= 1579409630;
assign addr[4787]= 1630224009;
assign addr[4788]= 1678970324;
assign addr[4789]= 1725586737;
assign addr[4790]= 1770014111;
assign addr[4791]= 1812196087;
assign addr[4792]= 1852079154;
assign addr[4793]= 1889612716;
assign addr[4794]= 1924749160;
assign addr[4795]= 1957443913;
assign addr[4796]= 1987655498;
assign addr[4797]= 2015345591;
assign addr[4798]= 2040479063;
assign addr[4799]= 2063024031;
assign addr[4800]= 2082951896;
assign addr[4801]= 2100237377;
assign addr[4802]= 2114858546;
assign addr[4803]= 2126796855;
assign addr[4804]= 2136037160;
assign addr[4805]= 2142567738;
assign addr[4806]= 2146380306;
assign addr[4807]= 2147470025;
assign addr[4808]= 2145835515;
assign addr[4809]= 2141478848;
assign addr[4810]= 2134405552;
assign addr[4811]= 2124624598;
assign addr[4812]= 2112148396;
assign addr[4813]= 2096992772;
assign addr[4814]= 2079176953;
assign addr[4815]= 2058723538;
assign addr[4816]= 2035658475;
assign addr[4817]= 2010011024;
assign addr[4818]= 1981813720;
assign addr[4819]= 1951102334;
assign addr[4820]= 1917915825;
assign addr[4821]= 1882296293;
assign addr[4822]= 1844288924;
assign addr[4823]= 1803941934;
assign addr[4824]= 1761306505;
assign addr[4825]= 1716436725;
assign addr[4826]= 1669389513;
assign addr[4827]= 1620224553;
assign addr[4828]= 1569004214;
assign addr[4829]= 1515793473;
assign addr[4830]= 1460659832;
assign addr[4831]= 1403673233;
assign addr[4832]= 1344905966;
assign addr[4833]= 1284432584;
assign addr[4834]= 1222329801;
assign addr[4835]= 1158676398;
assign addr[4836]= 1093553126;
assign addr[4837]= 1027042599;
assign addr[4838]= 959229189;
assign addr[4839]= 890198924;
assign addr[4840]= 820039373;
assign addr[4841]= 748839539;
assign addr[4842]= 676689746;
assign addr[4843]= 603681519;
assign addr[4844]= 529907477;
assign addr[4845]= 455461206;
assign addr[4846]= 380437148;
assign addr[4847]= 304930476;
assign addr[4848]= 229036977;
assign addr[4849]= 152852926;
assign addr[4850]= 76474970;
assign addr[4851]= 0;
assign addr[4852]= -76474970;
assign addr[4853]= -152852926;
assign addr[4854]= -229036977;
assign addr[4855]= -304930476;
assign addr[4856]= -380437148;
assign addr[4857]= -455461206;
assign addr[4858]= -529907477;
assign addr[4859]= -603681519;
assign addr[4860]= -676689746;
assign addr[4861]= -748839539;
assign addr[4862]= -820039373;
assign addr[4863]= -890198924;
assign addr[4864]= -959229189;
assign addr[4865]= -1027042599;
assign addr[4866]= -1093553126;
assign addr[4867]= -1158676398;
assign addr[4868]= -1222329801;
assign addr[4869]= -1284432584;
assign addr[4870]= -1344905966;
assign addr[4871]= -1403673233;
assign addr[4872]= -1460659832;
assign addr[4873]= -1515793473;
assign addr[4874]= -1569004214;
assign addr[4875]= -1620224553;
assign addr[4876]= -1669389513;
assign addr[4877]= -1716436725;
assign addr[4878]= -1761306505;
assign addr[4879]= -1803941934;
assign addr[4880]= -1844288924;
assign addr[4881]= -1882296293;
assign addr[4882]= -1917915825;
assign addr[4883]= -1951102334;
assign addr[4884]= -1981813720;
assign addr[4885]= -2010011024;
assign addr[4886]= -2035658475;
assign addr[4887]= -2058723538;
assign addr[4888]= -2079176953;
assign addr[4889]= -2096992772;
assign addr[4890]= -2112148396;
assign addr[4891]= -2124624598;
assign addr[4892]= -2134405552;
assign addr[4893]= -2141478848;
assign addr[4894]= -2145835515;
assign addr[4895]= -2147470025;
assign addr[4896]= -2146380306;
assign addr[4897]= -2142567738;
assign addr[4898]= -2136037160;
assign addr[4899]= -2126796855;
assign addr[4900]= -2114858546;
assign addr[4901]= -2100237377;
assign addr[4902]= -2082951896;
assign addr[4903]= -2063024031;
assign addr[4904]= -2040479063;
assign addr[4905]= -2015345591;
assign addr[4906]= -1987655498;
assign addr[4907]= -1957443913;
assign addr[4908]= -1924749160;
assign addr[4909]= -1889612716;
assign addr[4910]= -1852079154;
assign addr[4911]= -1812196087;
assign addr[4912]= -1770014111;
assign addr[4913]= -1725586737;
assign addr[4914]= -1678970324;
assign addr[4915]= -1630224009;
assign addr[4916]= -1579409630;
assign addr[4917]= -1526591649;
assign addr[4918]= -1471837070;
assign addr[4919]= -1415215352;
assign addr[4920]= -1356798326;
assign addr[4921]= -1296660098;
assign addr[4922]= -1234876957;
assign addr[4923]= -1171527280;
assign addr[4924]= -1106691431;
assign addr[4925]= -1040451659;
assign addr[4926]= -972891995;
assign addr[4927]= -904098143;
assign addr[4928]= -834157373;
assign addr[4929]= -763158411;
assign addr[4930]= -691191324;
assign addr[4931]= -618347408;
assign addr[4932]= -544719071;
assign addr[4933]= -470399716;
assign addr[4934]= -395483624;
assign addr[4935]= -320065829;
assign addr[4936]= -244242007;
assign addr[4937]= -168108346;
assign addr[4938]= -91761426;
assign addr[4939]= -15298099;
assign addr[4940]= 61184634;
assign addr[4941]= 137589750;
assign addr[4942]= 213820322;
assign addr[4943]= 289779648;
assign addr[4944]= 365371365;
assign addr[4945]= 440499581;
assign addr[4946]= 515068990;
assign addr[4947]= 588984994;
assign addr[4948]= 662153826;
assign addr[4949]= 734482665;
assign addr[4950]= 805879757;
assign addr[4951]= 876254528;
assign addr[4952]= 945517704;
assign addr[4953]= 1013581418;
assign addr[4954]= 1080359326;
assign addr[4955]= 1145766716;
assign addr[4956]= 1209720613;
assign addr[4957]= 1272139887;
assign addr[4958]= 1332945355;
assign addr[4959]= 1392059879;
assign addr[4960]= 1449408469;
assign addr[4961]= 1504918373;
assign addr[4962]= 1558519173;
assign addr[4963]= 1610142873;
assign addr[4964]= 1659723983;
assign addr[4965]= 1707199606;
assign addr[4966]= 1752509516;
assign addr[4967]= 1795596234;
assign addr[4968]= 1836405100;
assign addr[4969]= 1874884346;
assign addr[4970]= 1910985158;
assign addr[4971]= 1944661739;
assign addr[4972]= 1975871368;
assign addr[4973]= 2004574453;
assign addr[4974]= 2030734582;
assign addr[4975]= 2054318569;
assign addr[4976]= 2075296495;
assign addr[4977]= 2093641749;
assign addr[4978]= 2109331059;
assign addr[4979]= 2122344521;
assign addr[4980]= 2132665626;
assign addr[4981]= 2140281282;
assign addr[4982]= 2145181827;
assign addr[4983]= 2147361045;
assign addr[4984]= 2146816171;
assign addr[4985]= 2143547897;
assign addr[4986]= 2137560369;
assign addr[4987]= 2128861181;
assign addr[4988]= 2117461370;
assign addr[4989]= 2103375398;
assign addr[4990]= 2086621133;
assign addr[4991]= 2067219829;
assign addr[4992]= 2045196100;
assign addr[4993]= 2020577882;
assign addr[4994]= 1993396407;
assign addr[4995]= 1963686155;
assign addr[4996]= 1931484818;
assign addr[4997]= 1896833245;
assign addr[4998]= 1859775393;
assign addr[4999]= 1820358275;
assign addr[5000]= 1778631892;
assign addr[5001]= 1734649179;
assign addr[5002]= 1688465931;
assign addr[5003]= 1640140734;
assign addr[5004]= 1589734894;
assign addr[5005]= 1537312353;
assign addr[5006]= 1482939614;
assign addr[5007]= 1426685652;
assign addr[5008]= 1368621831;
assign addr[5009]= 1308821808;
assign addr[5010]= 1247361445;
assign addr[5011]= 1184318708;
assign addr[5012]= 1119773573;
assign addr[5013]= 1053807919;
assign addr[5014]= 986505429;
assign addr[5015]= 917951481;
assign addr[5016]= 848233042;
assign addr[5017]= 777438554;
assign addr[5018]= 705657826;
assign addr[5019]= 632981917;
assign addr[5020]= 559503022;
assign addr[5021]= 485314355;
assign addr[5022]= 410510029;
assign addr[5023]= 335184940;
assign addr[5024]= 259434643;
assign addr[5025]= 183355234;
assign addr[5026]= 107043224;
assign addr[5027]= 30595422;
assign addr[5028]= -45891193;
assign addr[5029]= -122319591;
assign addr[5030]= -198592817;
assign addr[5031]= -274614114;
assign addr[5032]= -350287041;
assign addr[5033]= -425515602;
assign addr[5034]= -500204365;
assign addr[5035]= -574258580;
assign addr[5036]= -647584304;
assign addr[5037]= -720088517;
assign addr[5038]= -791679244;
assign addr[5039]= -862265664;
assign addr[5040]= -931758235;
assign addr[5041]= -1000068799;
assign addr[5042]= -1067110699;
assign addr[5043]= -1132798888;
assign addr[5044]= -1197050035;
assign addr[5045]= -1259782632;
assign addr[5046]= -1320917099;
assign addr[5047]= -1380375881;
assign addr[5048]= -1438083551;
assign addr[5049]= -1493966902;
assign addr[5050]= -1547955041;
assign addr[5051]= -1599979481;
assign addr[5052]= -1649974225;
assign addr[5053]= -1697875851;
assign addr[5054]= -1743623590;
assign addr[5055]= -1787159411;
assign addr[5056]= -1828428082;
assign addr[5057]= -1867377253;
assign addr[5058]= -1903957513;
assign addr[5059]= -1938122457;
assign addr[5060]= -1969828744;
assign addr[5061]= -1999036154;
assign addr[5062]= -2025707632;
assign addr[5063]= -2049809346;
assign addr[5064]= -2071310720;
assign addr[5065]= -2090184478;
assign addr[5066]= -2106406677;
assign addr[5067]= -2119956737;
assign addr[5068]= -2130817471;
assign addr[5069]= -2138975100;
assign addr[5070]= -2144419275;
assign addr[5071]= -2147143090;
assign addr[5072]= -2147143090;
assign addr[5073]= -2144419275;
assign addr[5074]= -2138975100;
assign addr[5075]= -2130817471;
assign addr[5076]= -2119956737;
assign addr[5077]= -2106406677;
assign addr[5078]= -2090184478;
assign addr[5079]= -2071310720;
assign addr[5080]= -2049809346;
assign addr[5081]= -2025707632;
assign addr[5082]= -1999036154;
assign addr[5083]= -1969828744;
assign addr[5084]= -1938122457;
assign addr[5085]= -1903957513;
assign addr[5086]= -1867377253;
assign addr[5087]= -1828428082;
assign addr[5088]= -1787159411;
assign addr[5089]= -1743623590;
assign addr[5090]= -1697875851;
assign addr[5091]= -1649974225;
assign addr[5092]= -1599979481;
assign addr[5093]= -1547955041;
assign addr[5094]= -1493966902;
assign addr[5095]= -1438083551;
assign addr[5096]= -1380375881;
assign addr[5097]= -1320917099;
assign addr[5098]= -1259782632;
assign addr[5099]= -1197050035;
assign addr[5100]= -1132798888;
assign addr[5101]= -1067110699;
assign addr[5102]= -1000068799;
assign addr[5103]= -931758235;
assign addr[5104]= -862265664;
assign addr[5105]= -791679244;
assign addr[5106]= -720088517;
assign addr[5107]= -647584304;
assign addr[5108]= -574258580;
assign addr[5109]= -500204365;
assign addr[5110]= -425515602;
assign addr[5111]= -350287041;
assign addr[5112]= -274614114;
assign addr[5113]= -198592817;
assign addr[5114]= -122319591;
assign addr[5115]= -45891193;
assign addr[5116]= 30595422;
assign addr[5117]= 107043224;
assign addr[5118]= 183355234;
assign addr[5119]= 259434643;
assign addr[5120]= 335184940;
assign addr[5121]= 410510029;
assign addr[5122]= 485314355;
assign addr[5123]= 559503022;
assign addr[5124]= 632981917;
assign addr[5125]= 705657826;
assign addr[5126]= 777438554;
assign addr[5127]= 848233042;
assign addr[5128]= 917951481;
assign addr[5129]= 986505429;
assign addr[5130]= 1053807919;
assign addr[5131]= 1119773573;
assign addr[5132]= 1184318708;
assign addr[5133]= 1247361445;
assign addr[5134]= 1308821808;
assign addr[5135]= 1368621831;
assign addr[5136]= 1426685652;
assign addr[5137]= 1482939614;
assign addr[5138]= 1537312353;
assign addr[5139]= 1589734894;
assign addr[5140]= 1640140734;
assign addr[5141]= 1688465931;
assign addr[5142]= 1734649179;
assign addr[5143]= 1778631892;
assign addr[5144]= 1820358275;
assign addr[5145]= 1859775393;
assign addr[5146]= 1896833245;
assign addr[5147]= 1931484818;
assign addr[5148]= 1963686155;
assign addr[5149]= 1993396407;
assign addr[5150]= 2020577882;
assign addr[5151]= 2045196100;
assign addr[5152]= 2067219829;
assign addr[5153]= 2086621133;
assign addr[5154]= 2103375398;
assign addr[5155]= 2117461370;
assign addr[5156]= 2128861181;
assign addr[5157]= 2137560369;
assign addr[5158]= 2143547897;
assign addr[5159]= 2146816171;
assign addr[5160]= 2147361045;
assign addr[5161]= 2145181827;
assign addr[5162]= 2140281282;
assign addr[5163]= 2132665626;
assign addr[5164]= 2122344521;
assign addr[5165]= 2109331059;
assign addr[5166]= 2093641749;
assign addr[5167]= 2075296495;
assign addr[5168]= 2054318569;
assign addr[5169]= 2030734582;
assign addr[5170]= 2004574453;
assign addr[5171]= 1975871368;
assign addr[5172]= 1944661739;
assign addr[5173]= 1910985158;
assign addr[5174]= 1874884346;
assign addr[5175]= 1836405100;
assign addr[5176]= 1795596234;
assign addr[5177]= 1752509516;
assign addr[5178]= 1707199606;
assign addr[5179]= 1659723983;
assign addr[5180]= 1610142873;
assign addr[5181]= 1558519173;
assign addr[5182]= 1504918373;
assign addr[5183]= 1449408469;
assign addr[5184]= 1392059879;
assign addr[5185]= 1332945355;
assign addr[5186]= 1272139887;
assign addr[5187]= 1209720613;
assign addr[5188]= 1145766716;
assign addr[5189]= 1080359326;
assign addr[5190]= 1013581418;
assign addr[5191]= 945517704;
assign addr[5192]= 876254528;
assign addr[5193]= 805879757;
assign addr[5194]= 734482665;
assign addr[5195]= 662153826;
assign addr[5196]= 588984994;
assign addr[5197]= 515068990;
assign addr[5198]= 440499581;
assign addr[5199]= 365371365;
assign addr[5200]= 289779648;
assign addr[5201]= 213820322;
assign addr[5202]= 137589750;
assign addr[5203]= 61184634;
assign addr[5204]= -15298099;
assign addr[5205]= -91761426;
assign addr[5206]= -168108346;
assign addr[5207]= -244242007;
assign addr[5208]= -320065829;
assign addr[5209]= -395483624;
assign addr[5210]= -470399716;
assign addr[5211]= -544719071;
assign addr[5212]= -618347408;
assign addr[5213]= -691191324;
assign addr[5214]= -763158411;
assign addr[5215]= -834157373;
assign addr[5216]= -904098143;
assign addr[5217]= -972891995;
assign addr[5218]= -1040451659;
assign addr[5219]= -1106691431;
assign addr[5220]= -1171527280;
assign addr[5221]= -1234876957;
assign addr[5222]= -1296660098;
assign addr[5223]= -1356798326;
assign addr[5224]= -1415215352;
assign addr[5225]= -1471837070;
assign addr[5226]= -1526591649;
assign addr[5227]= -1579409630;
assign addr[5228]= -1630224009;
assign addr[5229]= -1678970324;
assign addr[5230]= -1725586737;
assign addr[5231]= -1770014111;
assign addr[5232]= -1812196087;
assign addr[5233]= -1852079154;
assign addr[5234]= -1889612716;
assign addr[5235]= -1924749160;
assign addr[5236]= -1957443913;
assign addr[5237]= -1987655498;
assign addr[5238]= -2015345591;
assign addr[5239]= -2040479063;
assign addr[5240]= -2063024031;
assign addr[5241]= -2082951896;
assign addr[5242]= -2100237377;
assign addr[5243]= -2114858546;
assign addr[5244]= -2126796855;
assign addr[5245]= -2136037160;
assign addr[5246]= -2142567738;
assign addr[5247]= -2146380306;
assign addr[5248]= -2147470025;
assign addr[5249]= -2145835515;
assign addr[5250]= -2141478848;
assign addr[5251]= -2134405552;
assign addr[5252]= -2124624598;
assign addr[5253]= -2112148396;
assign addr[5254]= -2096992772;
assign addr[5255]= -2079176953;
assign addr[5256]= -2058723538;
assign addr[5257]= -2035658475;
assign addr[5258]= -2010011024;
assign addr[5259]= -1981813720;
assign addr[5260]= -1951102334;
assign addr[5261]= -1917915825;
assign addr[5262]= -1882296293;
assign addr[5263]= -1844288924;
assign addr[5264]= -1803941934;
assign addr[5265]= -1761306505;
assign addr[5266]= -1716436725;
assign addr[5267]= -1669389513;
assign addr[5268]= -1620224553;
assign addr[5269]= -1569004214;
assign addr[5270]= -1515793473;
assign addr[5271]= -1460659832;
assign addr[5272]= -1403673233;
assign addr[5273]= -1344905966;
assign addr[5274]= -1284432584;
assign addr[5275]= -1222329801;
assign addr[5276]= -1158676398;
assign addr[5277]= -1093553126;
assign addr[5278]= -1027042599;
assign addr[5279]= -959229189;
assign addr[5280]= -890198924;
assign addr[5281]= -820039373;
assign addr[5282]= -748839539;
assign addr[5283]= -676689746;
assign addr[5284]= -603681519;
assign addr[5285]= -529907477;
assign addr[5286]= -455461206;
assign addr[5287]= -380437148;
assign addr[5288]= -304930476;
assign addr[5289]= -229036977;
assign addr[5290]= -152852926;
assign addr[5291]= -76474970;
assign addr[5292]= 0;
assign addr[5293]= 76474970;
assign addr[5294]= 152852926;
assign addr[5295]= 229036977;
assign addr[5296]= 304930476;
assign addr[5297]= 380437148;
assign addr[5298]= 455461206;
assign addr[5299]= 529907477;
assign addr[5300]= 603681519;
assign addr[5301]= 676689746;
assign addr[5302]= 748839539;
assign addr[5303]= 820039373;
assign addr[5304]= 890198924;
assign addr[5305]= 959229189;
assign addr[5306]= 1027042599;
assign addr[5307]= 1093553126;
assign addr[5308]= 1158676398;
assign addr[5309]= 1222329801;
assign addr[5310]= 1284432584;
assign addr[5311]= 1344905966;
assign addr[5312]= 1403673233;
assign addr[5313]= 1460659832;
assign addr[5314]= 1515793473;
assign addr[5315]= 1569004214;
assign addr[5316]= 1620224553;
assign addr[5317]= 1669389513;
assign addr[5318]= 1716436725;
assign addr[5319]= 1761306505;
assign addr[5320]= 1803941934;
assign addr[5321]= 1844288924;
assign addr[5322]= 1882296293;
assign addr[5323]= 1917915825;
assign addr[5324]= 1951102334;
assign addr[5325]= 1981813720;
assign addr[5326]= 2010011024;
assign addr[5327]= 2035658475;
assign addr[5328]= 2058723538;
assign addr[5329]= 2079176953;
assign addr[5330]= 2096992772;
assign addr[5331]= 2112148396;
assign addr[5332]= 2124624598;
assign addr[5333]= 2134405552;
assign addr[5334]= 2141478848;
assign addr[5335]= 2145835515;
assign addr[5336]= 2147470025;
assign addr[5337]= 2146380306;
assign addr[5338]= 2142567738;
assign addr[5339]= 2136037160;
assign addr[5340]= 2126796855;
assign addr[5341]= 2114858546;
assign addr[5342]= 2100237377;
assign addr[5343]= 2082951896;
assign addr[5344]= 2063024031;
assign addr[5345]= 2040479063;
assign addr[5346]= 2015345591;
assign addr[5347]= 1987655498;
assign addr[5348]= 1957443913;
assign addr[5349]= 1924749160;
assign addr[5350]= 1889612716;
assign addr[5351]= 1852079154;
assign addr[5352]= 1812196087;
assign addr[5353]= 1770014111;
assign addr[5354]= 1725586737;
assign addr[5355]= 1678970324;
assign addr[5356]= 1630224009;
assign addr[5357]= 1579409630;
assign addr[5358]= 1526591649;
assign addr[5359]= 1471837070;
assign addr[5360]= 1415215352;
assign addr[5361]= 1356798326;
assign addr[5362]= 1296660098;
assign addr[5363]= 1234876957;
assign addr[5364]= 1171527280;
assign addr[5365]= 1106691431;
assign addr[5366]= 1040451659;
assign addr[5367]= 972891995;
assign addr[5368]= 904098143;
assign addr[5369]= 834157373;
assign addr[5370]= 763158411;
assign addr[5371]= 691191324;
assign addr[5372]= 618347408;
assign addr[5373]= 544719071;
assign addr[5374]= 470399716;
assign addr[5375]= 395483624;
assign addr[5376]= 320065829;
assign addr[5377]= 244242007;
assign addr[5378]= 168108346;
assign addr[5379]= 91761426;
assign addr[5380]= 15298099;
assign addr[5381]= -61184634;
assign addr[5382]= -137589750;
assign addr[5383]= -213820322;
assign addr[5384]= -289779648;
assign addr[5385]= -365371365;
assign addr[5386]= -440499581;
assign addr[5387]= -515068990;
assign addr[5388]= -588984994;
assign addr[5389]= -662153826;
assign addr[5390]= -734482665;
assign addr[5391]= -805879757;
assign addr[5392]= -876254528;
assign addr[5393]= -945517704;
assign addr[5394]= -1013581418;
assign addr[5395]= -1080359326;
assign addr[5396]= -1145766716;
assign addr[5397]= -1209720613;
assign addr[5398]= -1272139887;
assign addr[5399]= -1332945355;
assign addr[5400]= -1392059879;
assign addr[5401]= -1449408469;
assign addr[5402]= -1504918373;
assign addr[5403]= -1558519173;
assign addr[5404]= -1610142873;
assign addr[5405]= -1659723983;
assign addr[5406]= -1707199606;
assign addr[5407]= -1752509516;
assign addr[5408]= -1795596234;
assign addr[5409]= -1836405100;
assign addr[5410]= -1874884346;
assign addr[5411]= -1910985158;
assign addr[5412]= -1944661739;
assign addr[5413]= -1975871368;
assign addr[5414]= -2004574453;
assign addr[5415]= -2030734582;
assign addr[5416]= -2054318569;
assign addr[5417]= -2075296495;
assign addr[5418]= -2093641749;
assign addr[5419]= -2109331059;
assign addr[5420]= -2122344521;
assign addr[5421]= -2132665626;
assign addr[5422]= -2140281282;
assign addr[5423]= -2145181827;
assign addr[5424]= -2147361045;
assign addr[5425]= -2146816171;
assign addr[5426]= -2143547897;
assign addr[5427]= -2137560369;
assign addr[5428]= -2128861181;
assign addr[5429]= -2117461370;
assign addr[5430]= -2103375398;
assign addr[5431]= -2086621133;
assign addr[5432]= -2067219829;
assign addr[5433]= -2045196100;
assign addr[5434]= -2020577882;
assign addr[5435]= -1993396407;
assign addr[5436]= -1963686155;
assign addr[5437]= -1931484818;
assign addr[5438]= -1896833245;
assign addr[5439]= -1859775393;
assign addr[5440]= -1820358275;
assign addr[5441]= -1778631892;
assign addr[5442]= -1734649179;
assign addr[5443]= -1688465931;
assign addr[5444]= -1640140734;
assign addr[5445]= -1589734894;
assign addr[5446]= -1537312353;
assign addr[5447]= -1482939614;
assign addr[5448]= -1426685652;
assign addr[5449]= -1368621831;
assign addr[5450]= -1308821808;
assign addr[5451]= -1247361445;
assign addr[5452]= -1184318708;
assign addr[5453]= -1119773573;
assign addr[5454]= -1053807919;
assign addr[5455]= -986505429;
assign addr[5456]= -917951481;
assign addr[5457]= -848233042;
assign addr[5458]= -777438554;
assign addr[5459]= -705657826;
assign addr[5460]= -632981917;
assign addr[5461]= -559503022;
assign addr[5462]= -485314355;
assign addr[5463]= -410510029;
assign addr[5464]= -335184940;
assign addr[5465]= -259434643;
assign addr[5466]= -183355234;
assign addr[5467]= -107043224;
assign addr[5468]= -30595422;
assign addr[5469]= 45891193;
assign addr[5470]= 122319591;
assign addr[5471]= 198592817;
assign addr[5472]= 274614114;
assign addr[5473]= 350287041;
assign addr[5474]= 425515602;
assign addr[5475]= 500204365;
assign addr[5476]= 574258580;
assign addr[5477]= 647584304;
assign addr[5478]= 720088517;
assign addr[5479]= 791679244;
assign addr[5480]= 862265664;
assign addr[5481]= 931758235;
assign addr[5482]= 1000068799;
assign addr[5483]= 1067110699;
assign addr[5484]= 1132798888;
assign addr[5485]= 1197050035;
assign addr[5486]= 1259782632;
assign addr[5487]= 1320917099;
assign addr[5488]= 1380375881;
assign addr[5489]= 1438083551;
assign addr[5490]= 1493966902;
assign addr[5491]= 1547955041;
assign addr[5492]= 1599979481;
assign addr[5493]= 1649974225;
assign addr[5494]= 1697875851;
assign addr[5495]= 1743623590;
assign addr[5496]= 1787159411;
assign addr[5497]= 1828428082;
assign addr[5498]= 1867377253;
assign addr[5499]= 1903957513;
assign addr[5500]= 1938122457;
assign addr[5501]= 1969828744;
assign addr[5502]= 1999036154;
assign addr[5503]= 2025707632;
assign addr[5504]= 2049809346;
assign addr[5505]= 2071310720;
assign addr[5506]= 2090184478;
assign addr[5507]= 2106406677;
assign addr[5508]= 2119956737;
assign addr[5509]= 2130817471;
assign addr[5510]= 2138975100;
assign addr[5511]= 2144419275;
assign addr[5512]= 2147143090;
assign addr[5513]= 2147143090;
assign addr[5514]= 2144419275;
assign addr[5515]= 2138975100;
assign addr[5516]= 2130817471;
assign addr[5517]= 2119956737;
assign addr[5518]= 2106406677;
assign addr[5519]= 2090184478;
assign addr[5520]= 2071310720;
assign addr[5521]= 2049809346;
assign addr[5522]= 2025707632;
assign addr[5523]= 1999036154;
assign addr[5524]= 1969828744;
assign addr[5525]= 1938122457;
assign addr[5526]= 1903957513;
assign addr[5527]= 1867377253;
assign addr[5528]= 1828428082;
assign addr[5529]= 1787159411;
assign addr[5530]= 1743623590;
assign addr[5531]= 1697875851;
assign addr[5532]= 1649974225;
assign addr[5533]= 1599979481;
assign addr[5534]= 1547955041;
assign addr[5535]= 1493966902;
assign addr[5536]= 1438083551;
assign addr[5537]= 1380375881;
assign addr[5538]= 1320917099;
assign addr[5539]= 1259782632;
assign addr[5540]= 1197050035;
assign addr[5541]= 1132798888;
assign addr[5542]= 1067110699;
assign addr[5543]= 1000068799;
assign addr[5544]= 931758235;
assign addr[5545]= 862265664;
assign addr[5546]= 791679244;
assign addr[5547]= 720088517;
assign addr[5548]= 647584304;
assign addr[5549]= 574258580;
assign addr[5550]= 500204365;
assign addr[5551]= 425515602;
assign addr[5552]= 350287041;
assign addr[5553]= 274614114;
assign addr[5554]= 198592817;
assign addr[5555]= 122319591;
assign addr[5556]= 45891193;
assign addr[5557]= -30595422;
assign addr[5558]= -107043224;
assign addr[5559]= -183355234;
assign addr[5560]= -259434643;
assign addr[5561]= -335184940;
assign addr[5562]= -410510029;
assign addr[5563]= -485314355;
assign addr[5564]= -559503022;
assign addr[5565]= -632981917;
assign addr[5566]= -705657826;
assign addr[5567]= -777438554;
assign addr[5568]= -848233042;
assign addr[5569]= -917951481;
assign addr[5570]= -986505429;
assign addr[5571]= -1053807919;
assign addr[5572]= -1119773573;
assign addr[5573]= -1184318708;
assign addr[5574]= -1247361445;
assign addr[5575]= -1308821808;
assign addr[5576]= -1368621831;
assign addr[5577]= -1426685652;
assign addr[5578]= -1482939614;
assign addr[5579]= -1537312353;
assign addr[5580]= -1589734894;
assign addr[5581]= -1640140734;
assign addr[5582]= -1688465931;
assign addr[5583]= -1734649179;
assign addr[5584]= -1778631892;
assign addr[5585]= -1820358275;
assign addr[5586]= -1859775393;
assign addr[5587]= -1896833245;
assign addr[5588]= -1931484818;
assign addr[5589]= -1963686155;
assign addr[5590]= -1993396407;
assign addr[5591]= -2020577882;
assign addr[5592]= -2045196100;
assign addr[5593]= -2067219829;
assign addr[5594]= -2086621133;
assign addr[5595]= -2103375398;
assign addr[5596]= -2117461370;
assign addr[5597]= -2128861181;
assign addr[5598]= -2137560369;
assign addr[5599]= -2143547897;
assign addr[5600]= -2146816171;
assign addr[5601]= -2147361045;
assign addr[5602]= -2145181827;
assign addr[5603]= -2140281282;
assign addr[5604]= -2132665626;
assign addr[5605]= -2122344521;
assign addr[5606]= -2109331059;
assign addr[5607]= -2093641749;
assign addr[5608]= -2075296495;
assign addr[5609]= -2054318569;
assign addr[5610]= -2030734582;
assign addr[5611]= -2004574453;
assign addr[5612]= -1975871368;
assign addr[5613]= -1944661739;
assign addr[5614]= -1910985158;
assign addr[5615]= -1874884346;
assign addr[5616]= -1836405100;
assign addr[5617]= -1795596234;
assign addr[5618]= -1752509516;
assign addr[5619]= -1707199606;
assign addr[5620]= -1659723983;
assign addr[5621]= -1610142873;
assign addr[5622]= -1558519173;
assign addr[5623]= -1504918373;
assign addr[5624]= -1449408469;
assign addr[5625]= -1392059879;
assign addr[5626]= -1332945355;
assign addr[5627]= -1272139887;
assign addr[5628]= -1209720613;
assign addr[5629]= -1145766716;
assign addr[5630]= -1080359326;
assign addr[5631]= -1013581418;
assign addr[5632]= -945517704;
assign addr[5633]= -876254528;
assign addr[5634]= -805879757;
assign addr[5635]= -734482665;
assign addr[5636]= -662153826;
assign addr[5637]= -588984994;
assign addr[5638]= -515068990;
assign addr[5639]= -440499581;
assign addr[5640]= -365371365;
assign addr[5641]= -289779648;
assign addr[5642]= -213820322;
assign addr[5643]= -137589750;
assign addr[5644]= -61184634;
assign addr[5645]= 15298099;
assign addr[5646]= 91761426;
assign addr[5647]= 168108346;
assign addr[5648]= 244242007;
assign addr[5649]= 320065829;
assign addr[5650]= 395483624;
assign addr[5651]= 470399716;
assign addr[5652]= 544719071;
assign addr[5653]= 618347408;
assign addr[5654]= 691191324;
assign addr[5655]= 763158411;
assign addr[5656]= 834157373;
assign addr[5657]= 904098143;
assign addr[5658]= 972891995;
assign addr[5659]= 1040451659;
assign addr[5660]= 1106691431;
assign addr[5661]= 1171527280;
assign addr[5662]= 1234876957;
assign addr[5663]= 1296660098;
assign addr[5664]= 1356798326;
assign addr[5665]= 1415215352;
assign addr[5666]= 1471837070;
assign addr[5667]= 1526591649;
assign addr[5668]= 1579409630;
assign addr[5669]= 1630224009;
assign addr[5670]= 1678970324;
assign addr[5671]= 1725586737;
assign addr[5672]= 1770014111;
assign addr[5673]= 1812196087;
assign addr[5674]= 1852079154;
assign addr[5675]= 1889612716;
assign addr[5676]= 1924749160;
assign addr[5677]= 1957443913;
assign addr[5678]= 1987655498;
assign addr[5679]= 2015345591;
assign addr[5680]= 2040479063;
assign addr[5681]= 2063024031;
assign addr[5682]= 2082951896;
assign addr[5683]= 2100237377;
assign addr[5684]= 2114858546;
assign addr[5685]= 2126796855;
assign addr[5686]= 2136037160;
assign addr[5687]= 2142567738;
assign addr[5688]= 2146380306;
assign addr[5689]= 2147470025;
assign addr[5690]= 2145835515;
assign addr[5691]= 2141478848;
assign addr[5692]= 2134405552;
assign addr[5693]= 2124624598;
assign addr[5694]= 2112148396;
assign addr[5695]= 2096992772;
assign addr[5696]= 2079176953;
assign addr[5697]= 2058723538;
assign addr[5698]= 2035658475;
assign addr[5699]= 2010011024;
assign addr[5700]= 1981813720;
assign addr[5701]= 1951102334;
assign addr[5702]= 1917915825;
assign addr[5703]= 1882296293;
assign addr[5704]= 1844288924;
assign addr[5705]= 1803941934;
assign addr[5706]= 1761306505;
assign addr[5707]= 1716436725;
assign addr[5708]= 1669389513;
assign addr[5709]= 1620224553;
assign addr[5710]= 1569004214;
assign addr[5711]= 1515793473;
assign addr[5712]= 1460659832;
assign addr[5713]= 1403673233;
assign addr[5714]= 1344905966;
assign addr[5715]= 1284432584;
assign addr[5716]= 1222329801;
assign addr[5717]= 1158676398;
assign addr[5718]= 1093553126;
assign addr[5719]= 1027042599;
assign addr[5720]= 959229189;
assign addr[5721]= 890198924;
assign addr[5722]= 820039373;
assign addr[5723]= 748839539;
assign addr[5724]= 676689746;
assign addr[5725]= 603681519;
assign addr[5726]= 529907477;
assign addr[5727]= 455461206;
assign addr[5728]= 380437148;
assign addr[5729]= 304930476;
assign addr[5730]= 229036977;
assign addr[5731]= 152852926;
assign addr[5732]= 76474970;
assign addr[5733]= 0;
assign addr[5734]= -76474970;
assign addr[5735]= -152852926;
assign addr[5736]= -229036977;
assign addr[5737]= -304930476;
assign addr[5738]= -380437148;
assign addr[5739]= -455461206;
assign addr[5740]= -529907477;
assign addr[5741]= -603681519;
assign addr[5742]= -676689746;
assign addr[5743]= -748839539;
assign addr[5744]= -820039373;
assign addr[5745]= -890198924;
assign addr[5746]= -959229189;
assign addr[5747]= -1027042599;
assign addr[5748]= -1093553126;
assign addr[5749]= -1158676398;
assign addr[5750]= -1222329801;
assign addr[5751]= -1284432584;
assign addr[5752]= -1344905966;
assign addr[5753]= -1403673233;
assign addr[5754]= -1460659832;
assign addr[5755]= -1515793473;
assign addr[5756]= -1569004214;
assign addr[5757]= -1620224553;
assign addr[5758]= -1669389513;
assign addr[5759]= -1716436725;
assign addr[5760]= -1761306505;
assign addr[5761]= -1803941934;
assign addr[5762]= -1844288924;
assign addr[5763]= -1882296293;
assign addr[5764]= -1917915825;
assign addr[5765]= -1951102334;
assign addr[5766]= -1981813720;
assign addr[5767]= -2010011024;
assign addr[5768]= -2035658475;
assign addr[5769]= -2058723538;
assign addr[5770]= -2079176953;
assign addr[5771]= -2096992772;
assign addr[5772]= -2112148396;
assign addr[5773]= -2124624598;
assign addr[5774]= -2134405552;
assign addr[5775]= -2141478848;
assign addr[5776]= -2145835515;
assign addr[5777]= -2147470025;
assign addr[5778]= -2146380306;
assign addr[5779]= -2142567738;
assign addr[5780]= -2136037160;
assign addr[5781]= -2126796855;
assign addr[5782]= -2114858546;
assign addr[5783]= -2100237377;
assign addr[5784]= -2082951896;
assign addr[5785]= -2063024031;
assign addr[5786]= -2040479063;
assign addr[5787]= -2015345591;
assign addr[5788]= -1987655498;
assign addr[5789]= -1957443913;
assign addr[5790]= -1924749160;
assign addr[5791]= -1889612716;
assign addr[5792]= -1852079154;
assign addr[5793]= -1812196087;
assign addr[5794]= -1770014111;
assign addr[5795]= -1725586737;
assign addr[5796]= -1678970324;
assign addr[5797]= -1630224009;
assign addr[5798]= -1579409630;
assign addr[5799]= -1526591649;
assign addr[5800]= -1471837070;
assign addr[5801]= -1415215352;
assign addr[5802]= -1356798326;
assign addr[5803]= -1296660098;
assign addr[5804]= -1234876957;
assign addr[5805]= -1171527280;
assign addr[5806]= -1106691431;
assign addr[5807]= -1040451659;
assign addr[5808]= -972891995;
assign addr[5809]= -904098143;
assign addr[5810]= -834157373;
assign addr[5811]= -763158411;
assign addr[5812]= -691191324;
assign addr[5813]= -618347408;
assign addr[5814]= -544719071;
assign addr[5815]= -470399716;
assign addr[5816]= -395483624;
assign addr[5817]= -320065829;
assign addr[5818]= -244242007;
assign addr[5819]= -168108346;
assign addr[5820]= -91761426;
assign addr[5821]= -15298099;
assign addr[5822]= 61184634;
assign addr[5823]= 137589750;
assign addr[5824]= 213820322;
assign addr[5825]= 289779648;
assign addr[5826]= 365371365;
assign addr[5827]= 440499581;
assign addr[5828]= 515068990;
assign addr[5829]= 588984994;
assign addr[5830]= 662153826;
assign addr[5831]= 734482665;
assign addr[5832]= 805879757;
assign addr[5833]= 876254528;
assign addr[5834]= 945517704;
assign addr[5835]= 1013581418;
assign addr[5836]= 1080359326;
assign addr[5837]= 1145766716;
assign addr[5838]= 1209720613;
assign addr[5839]= 1272139887;
assign addr[5840]= 1332945355;
assign addr[5841]= 1392059879;
assign addr[5842]= 1449408469;
assign addr[5843]= 1504918373;
assign addr[5844]= 1558519173;
assign addr[5845]= 1610142873;
assign addr[5846]= 1659723983;
assign addr[5847]= 1707199606;
assign addr[5848]= 1752509516;
assign addr[5849]= 1795596234;
assign addr[5850]= 1836405100;
assign addr[5851]= 1874884346;
assign addr[5852]= 1910985158;
assign addr[5853]= 1944661739;
assign addr[5854]= 1975871368;
assign addr[5855]= 2004574453;
assign addr[5856]= 2030734582;
assign addr[5857]= 2054318569;
assign addr[5858]= 2075296495;
assign addr[5859]= 2093641749;
assign addr[5860]= 2109331059;
assign addr[5861]= 2122344521;
assign addr[5862]= 2132665626;
assign addr[5863]= 2140281282;
assign addr[5864]= 2145181827;
assign addr[5865]= 2147361045;
assign addr[5866]= 2146816171;
assign addr[5867]= 2143547897;
assign addr[5868]= 2137560369;
assign addr[5869]= 2128861181;
assign addr[5870]= 2117461370;
assign addr[5871]= 2103375398;
assign addr[5872]= 2086621133;
assign addr[5873]= 2067219829;
assign addr[5874]= 2045196100;
assign addr[5875]= 2020577882;
assign addr[5876]= 1993396407;
assign addr[5877]= 1963686155;
assign addr[5878]= 1931484818;
assign addr[5879]= 1896833245;
assign addr[5880]= 1859775393;
assign addr[5881]= 1820358275;
assign addr[5882]= 1778631892;
assign addr[5883]= 1734649179;
assign addr[5884]= 1688465931;
assign addr[5885]= 1640140734;
assign addr[5886]= 1589734894;
assign addr[5887]= 1537312353;
assign addr[5888]= 1482939614;
assign addr[5889]= 1426685652;
assign addr[5890]= 1368621831;
assign addr[5891]= 1308821808;
assign addr[5892]= 1247361445;
assign addr[5893]= 1184318708;
assign addr[5894]= 1119773573;
assign addr[5895]= 1053807919;
assign addr[5896]= 986505429;
assign addr[5897]= 917951481;
assign addr[5898]= 848233042;
assign addr[5899]= 777438554;
assign addr[5900]= 705657826;
assign addr[5901]= 632981917;
assign addr[5902]= 559503022;
assign addr[5903]= 485314355;
assign addr[5904]= 410510029;
assign addr[5905]= 335184940;
assign addr[5906]= 259434643;
assign addr[5907]= 183355234;
assign addr[5908]= 107043224;
assign addr[5909]= 30595422;
assign addr[5910]= -45891193;
assign addr[5911]= -122319591;
assign addr[5912]= -198592817;
assign addr[5913]= -274614114;
assign addr[5914]= -350287041;
assign addr[5915]= -425515602;
assign addr[5916]= -500204365;
assign addr[5917]= -574258580;
assign addr[5918]= -647584304;
assign addr[5919]= -720088517;
assign addr[5920]= -791679244;
assign addr[5921]= -862265664;
assign addr[5922]= -931758235;
assign addr[5923]= -1000068799;
assign addr[5924]= -1067110699;
assign addr[5925]= -1132798888;
assign addr[5926]= -1197050035;
assign addr[5927]= -1259782632;
assign addr[5928]= -1320917099;
assign addr[5929]= -1380375881;
assign addr[5930]= -1438083551;
assign addr[5931]= -1493966902;
assign addr[5932]= -1547955041;
assign addr[5933]= -1599979481;
assign addr[5934]= -1649974225;
assign addr[5935]= -1697875851;
assign addr[5936]= -1743623590;
assign addr[5937]= -1787159411;
assign addr[5938]= -1828428082;
assign addr[5939]= -1867377253;
assign addr[5940]= -1903957513;
assign addr[5941]= -1938122457;
assign addr[5942]= -1969828744;
assign addr[5943]= -1999036154;
assign addr[5944]= -2025707632;
assign addr[5945]= -2049809346;
assign addr[5946]= -2071310720;
assign addr[5947]= -2090184478;
assign addr[5948]= -2106406677;
assign addr[5949]= -2119956737;
assign addr[5950]= -2130817471;
assign addr[5951]= -2138975100;
assign addr[5952]= -2144419275;
assign addr[5953]= -2147143090;
assign addr[5954]= -2147143090;
assign addr[5955]= -2144419275;
assign addr[5956]= -2138975100;
assign addr[5957]= -2130817471;
assign addr[5958]= -2119956737;
assign addr[5959]= -2106406677;
assign addr[5960]= -2090184478;
assign addr[5961]= -2071310720;
assign addr[5962]= -2049809346;
assign addr[5963]= -2025707632;
assign addr[5964]= -1999036154;
assign addr[5965]= -1969828744;
assign addr[5966]= -1938122457;
assign addr[5967]= -1903957513;
assign addr[5968]= -1867377253;
assign addr[5969]= -1828428082;
assign addr[5970]= -1787159411;
assign addr[5971]= -1743623590;
assign addr[5972]= -1697875851;
assign addr[5973]= -1649974225;
assign addr[5974]= -1599979481;
assign addr[5975]= -1547955041;
assign addr[5976]= -1493966902;
assign addr[5977]= -1438083551;
assign addr[5978]= -1380375881;
assign addr[5979]= -1320917099;
assign addr[5980]= -1259782632;
assign addr[5981]= -1197050035;
assign addr[5982]= -1132798888;
assign addr[5983]= -1067110699;
assign addr[5984]= -1000068799;
assign addr[5985]= -931758235;
assign addr[5986]= -862265664;
assign addr[5987]= -791679244;
assign addr[5988]= -720088517;
assign addr[5989]= -647584304;
assign addr[5990]= -574258580;
assign addr[5991]= -500204365;
assign addr[5992]= -425515602;
assign addr[5993]= -350287041;
assign addr[5994]= -274614114;
assign addr[5995]= -198592817;
assign addr[5996]= -122319591;
assign addr[5997]= -45891193;
assign addr[5998]= 30595422;
assign addr[5999]= 107043224;
assign addr[6000]= 183355234;
assign addr[6001]= 259434643;
assign addr[6002]= 335184940;
assign addr[6003]= 410510029;
assign addr[6004]= 485314355;
assign addr[6005]= 559503022;
assign addr[6006]= 632981917;
assign addr[6007]= 705657826;
assign addr[6008]= 777438554;
assign addr[6009]= 848233042;
assign addr[6010]= 917951481;
assign addr[6011]= 986505429;
assign addr[6012]= 1053807919;
assign addr[6013]= 1119773573;
assign addr[6014]= 1184318708;
assign addr[6015]= 1247361445;
assign addr[6016]= 1308821808;
assign addr[6017]= 1368621831;
assign addr[6018]= 1426685652;
assign addr[6019]= 1482939614;
assign addr[6020]= 1537312353;
assign addr[6021]= 1589734894;
assign addr[6022]= 1640140734;
assign addr[6023]= 1688465931;
assign addr[6024]= 1734649179;
assign addr[6025]= 1778631892;
assign addr[6026]= 1820358275;
assign addr[6027]= 1859775393;
assign addr[6028]= 1896833245;
assign addr[6029]= 1931484818;
assign addr[6030]= 1963686155;
assign addr[6031]= 1993396407;
assign addr[6032]= 2020577882;
assign addr[6033]= 2045196100;
assign addr[6034]= 2067219829;
assign addr[6035]= 2086621133;
assign addr[6036]= 2103375398;
assign addr[6037]= 2117461370;
assign addr[6038]= 2128861181;
assign addr[6039]= 2137560369;
assign addr[6040]= 2143547897;
assign addr[6041]= 2146816171;
assign addr[6042]= 2147361045;
assign addr[6043]= 2145181827;
assign addr[6044]= 2140281282;
assign addr[6045]= 2132665626;
assign addr[6046]= 2122344521;
assign addr[6047]= 2109331059;
assign addr[6048]= 2093641749;
assign addr[6049]= 2075296495;
assign addr[6050]= 2054318569;
assign addr[6051]= 2030734582;
assign addr[6052]= 2004574453;
assign addr[6053]= 1975871368;
assign addr[6054]= 1944661739;
assign addr[6055]= 1910985158;
assign addr[6056]= 1874884346;
assign addr[6057]= 1836405100;
assign addr[6058]= 1795596234;
assign addr[6059]= 1752509516;
assign addr[6060]= 1707199606;
assign addr[6061]= 1659723983;
assign addr[6062]= 1610142873;
assign addr[6063]= 1558519173;
assign addr[6064]= 1504918373;
assign addr[6065]= 1449408469;
assign addr[6066]= 1392059879;
assign addr[6067]= 1332945355;
assign addr[6068]= 1272139887;
assign addr[6069]= 1209720613;
assign addr[6070]= 1145766716;
assign addr[6071]= 1080359326;
assign addr[6072]= 1013581418;
assign addr[6073]= 945517704;
assign addr[6074]= 876254528;
assign addr[6075]= 805879757;
assign addr[6076]= 734482665;
assign addr[6077]= 662153826;
assign addr[6078]= 588984994;
assign addr[6079]= 515068990;
assign addr[6080]= 440499581;
assign addr[6081]= 365371365;
assign addr[6082]= 289779648;
assign addr[6083]= 213820322;
assign addr[6084]= 137589750;
assign addr[6085]= 61184634;
assign addr[6086]= -15298099;
assign addr[6087]= -91761426;
assign addr[6088]= -168108346;
assign addr[6089]= -244242007;
assign addr[6090]= -320065829;
assign addr[6091]= -395483624;
assign addr[6092]= -470399716;
assign addr[6093]= -544719071;
assign addr[6094]= -618347408;
assign addr[6095]= -691191324;
assign addr[6096]= -763158411;
assign addr[6097]= -834157373;
assign addr[6098]= -904098143;
assign addr[6099]= -972891995;
assign addr[6100]= -1040451659;
assign addr[6101]= -1106691431;
assign addr[6102]= -1171527280;
assign addr[6103]= -1234876957;
assign addr[6104]= -1296660098;
assign addr[6105]= -1356798326;
assign addr[6106]= -1415215352;
assign addr[6107]= -1471837070;
assign addr[6108]= -1526591649;
assign addr[6109]= -1579409630;
assign addr[6110]= -1630224009;
assign addr[6111]= -1678970324;
assign addr[6112]= -1725586737;
assign addr[6113]= -1770014111;
assign addr[6114]= -1812196087;
assign addr[6115]= -1852079154;
assign addr[6116]= -1889612716;
assign addr[6117]= -1924749160;
assign addr[6118]= -1957443913;
assign addr[6119]= -1987655498;
assign addr[6120]= -2015345591;
assign addr[6121]= -2040479063;
assign addr[6122]= -2063024031;
assign addr[6123]= -2082951896;
assign addr[6124]= -2100237377;
assign addr[6125]= -2114858546;
assign addr[6126]= -2126796855;
assign addr[6127]= -2136037160;
assign addr[6128]= -2142567738;
assign addr[6129]= -2146380306;
assign addr[6130]= -2147470025;
assign addr[6131]= -2145835515;
assign addr[6132]= -2141478848;
assign addr[6133]= -2134405552;
assign addr[6134]= -2124624598;
assign addr[6135]= -2112148396;
assign addr[6136]= -2096992772;
assign addr[6137]= -2079176953;
assign addr[6138]= -2058723538;
assign addr[6139]= -2035658475;
assign addr[6140]= -2010011024;
assign addr[6141]= -1981813720;
assign addr[6142]= -1951102334;
assign addr[6143]= -1917915825;
assign addr[6144]= -1882296293;
assign addr[6145]= -1844288924;
assign addr[6146]= -1803941934;
assign addr[6147]= -1761306505;
assign addr[6148]= -1716436725;
assign addr[6149]= -1669389513;
assign addr[6150]= -1620224553;
assign addr[6151]= -1569004214;
assign addr[6152]= -1515793473;
assign addr[6153]= -1460659832;
assign addr[6154]= -1403673233;
assign addr[6155]= -1344905966;
assign addr[6156]= -1284432584;
assign addr[6157]= -1222329801;
assign addr[6158]= -1158676398;
assign addr[6159]= -1093553126;
assign addr[6160]= -1027042599;
assign addr[6161]= -959229189;
assign addr[6162]= -890198924;
assign addr[6163]= -820039373;
assign addr[6164]= -748839539;
assign addr[6165]= -676689746;
assign addr[6166]= -603681519;
assign addr[6167]= -529907477;
assign addr[6168]= -455461206;
assign addr[6169]= -380437148;
assign addr[6170]= -304930476;
assign addr[6171]= -229036977;
assign addr[6172]= -152852926;
assign addr[6173]= -76474970;
assign addr[6174]= 0;
assign addr[6175]= 76474970;
assign addr[6176]= 152852926;
assign addr[6177]= 229036977;
assign addr[6178]= 304930476;
assign addr[6179]= 380437148;
assign addr[6180]= 455461206;
assign addr[6181]= 529907477;
assign addr[6182]= 603681519;
assign addr[6183]= 676689746;
assign addr[6184]= 748839539;
assign addr[6185]= 820039373;
assign addr[6186]= 890198924;
assign addr[6187]= 959229189;
assign addr[6188]= 1027042599;
assign addr[6189]= 1093553126;
assign addr[6190]= 1158676398;
assign addr[6191]= 1222329801;
assign addr[6192]= 1284432584;
assign addr[6193]= 1344905966;
assign addr[6194]= 1403673233;
assign addr[6195]= 1460659832;
assign addr[6196]= 1515793473;
assign addr[6197]= 1569004214;
assign addr[6198]= 1620224553;
assign addr[6199]= 1669389513;
assign addr[6200]= 1716436725;
assign addr[6201]= 1761306505;
assign addr[6202]= 1803941934;
assign addr[6203]= 1844288924;
assign addr[6204]= 1882296293;
assign addr[6205]= 1917915825;
assign addr[6206]= 1951102334;
assign addr[6207]= 1981813720;
assign addr[6208]= 2010011024;
assign addr[6209]= 2035658475;
assign addr[6210]= 2058723538;
assign addr[6211]= 2079176953;
assign addr[6212]= 2096992772;
assign addr[6213]= 2112148396;
assign addr[6214]= 2124624598;
assign addr[6215]= 2134405552;
assign addr[6216]= 2141478848;
assign addr[6217]= 2145835515;
assign addr[6218]= 2147470025;
assign addr[6219]= 2146380306;
assign addr[6220]= 2142567738;
assign addr[6221]= 2136037160;
assign addr[6222]= 2126796855;
assign addr[6223]= 2114858546;
assign addr[6224]= 2100237377;
assign addr[6225]= 2082951896;
assign addr[6226]= 2063024031;
assign addr[6227]= 2040479063;
assign addr[6228]= 2015345591;
assign addr[6229]= 1987655498;
assign addr[6230]= 1957443913;
assign addr[6231]= 1924749160;
assign addr[6232]= 1889612716;
assign addr[6233]= 1852079154;
assign addr[6234]= 1812196087;
assign addr[6235]= 1770014111;
assign addr[6236]= 1725586737;
assign addr[6237]= 1678970324;
assign addr[6238]= 1630224009;
assign addr[6239]= 1579409630;
assign addr[6240]= 1526591649;
assign addr[6241]= 1471837070;
assign addr[6242]= 1415215352;
assign addr[6243]= 1356798326;
assign addr[6244]= 1296660098;
assign addr[6245]= 1234876957;
assign addr[6246]= 1171527280;
assign addr[6247]= 1106691431;
assign addr[6248]= 1040451659;
assign addr[6249]= 972891995;
assign addr[6250]= 904098143;
assign addr[6251]= 834157373;
assign addr[6252]= 763158411;
assign addr[6253]= 691191324;
assign addr[6254]= 618347408;
assign addr[6255]= 544719071;
assign addr[6256]= 470399716;
assign addr[6257]= 395483624;
assign addr[6258]= 320065829;
assign addr[6259]= 244242007;
assign addr[6260]= 168108346;
assign addr[6261]= 91761426;
assign addr[6262]= 15298099;
assign addr[6263]= -61184634;
assign addr[6264]= -137589750;
assign addr[6265]= -213820322;
assign addr[6266]= -289779648;
assign addr[6267]= -365371365;
assign addr[6268]= -440499581;
assign addr[6269]= -515068990;
assign addr[6270]= -588984994;
assign addr[6271]= -662153826;
assign addr[6272]= -734482665;
assign addr[6273]= -805879757;
assign addr[6274]= -876254528;
assign addr[6275]= -945517704;
assign addr[6276]= -1013581418;
assign addr[6277]= -1080359326;
assign addr[6278]= -1145766716;
assign addr[6279]= -1209720613;
assign addr[6280]= -1272139887;
assign addr[6281]= -1332945355;
assign addr[6282]= -1392059879;
assign addr[6283]= -1449408469;
assign addr[6284]= -1504918373;
assign addr[6285]= -1558519173;
assign addr[6286]= -1610142873;
assign addr[6287]= -1659723983;
assign addr[6288]= -1707199606;
assign addr[6289]= -1752509516;
assign addr[6290]= -1795596234;
assign addr[6291]= -1836405100;
assign addr[6292]= -1874884346;
assign addr[6293]= -1910985158;
assign addr[6294]= -1944661739;
assign addr[6295]= -1975871368;
assign addr[6296]= -2004574453;
assign addr[6297]= -2030734582;
assign addr[6298]= -2054318569;
assign addr[6299]= -2075296495;
assign addr[6300]= -2093641749;
assign addr[6301]= -2109331059;
assign addr[6302]= -2122344521;
assign addr[6303]= -2132665626;
assign addr[6304]= -2140281282;
assign addr[6305]= -2145181827;
assign addr[6306]= -2147361045;
assign addr[6307]= -2146816171;
assign addr[6308]= -2143547897;
assign addr[6309]= -2137560369;
assign addr[6310]= -2128861181;
assign addr[6311]= -2117461370;
assign addr[6312]= -2103375398;
assign addr[6313]= -2086621133;
assign addr[6314]= -2067219829;
assign addr[6315]= -2045196100;
assign addr[6316]= -2020577882;
assign addr[6317]= -1993396407;
assign addr[6318]= -1963686155;
assign addr[6319]= -1931484818;
assign addr[6320]= -1896833245;
assign addr[6321]= -1859775393;
assign addr[6322]= -1820358275;
assign addr[6323]= -1778631892;
assign addr[6324]= -1734649179;
assign addr[6325]= -1688465931;
assign addr[6326]= -1640140734;
assign addr[6327]= -1589734894;
assign addr[6328]= -1537312353;
assign addr[6329]= -1482939614;
assign addr[6330]= -1426685652;
assign addr[6331]= -1368621831;
assign addr[6332]= -1308821808;
assign addr[6333]= -1247361445;
assign addr[6334]= -1184318708;
assign addr[6335]= -1119773573;
assign addr[6336]= -1053807919;
assign addr[6337]= -986505429;
assign addr[6338]= -917951481;
assign addr[6339]= -848233042;
assign addr[6340]= -777438554;
assign addr[6341]= -705657826;
assign addr[6342]= -632981917;
assign addr[6343]= -559503022;
assign addr[6344]= -485314355;
assign addr[6345]= -410510029;
assign addr[6346]= -335184940;
assign addr[6347]= -259434643;
assign addr[6348]= -183355234;
assign addr[6349]= -107043224;
assign addr[6350]= -30595422;
assign addr[6351]= 45891193;
assign addr[6352]= 122319591;
assign addr[6353]= 198592817;
assign addr[6354]= 274614114;
assign addr[6355]= 350287041;
assign addr[6356]= 425515602;
assign addr[6357]= 500204365;
assign addr[6358]= 574258580;
assign addr[6359]= 647584304;
assign addr[6360]= 720088517;
assign addr[6361]= 791679244;
assign addr[6362]= 862265664;
assign addr[6363]= 931758235;
assign addr[6364]= 1000068799;
assign addr[6365]= 1067110699;
assign addr[6366]= 1132798888;
assign addr[6367]= 1197050035;
assign addr[6368]= 1259782632;
assign addr[6369]= 1320917099;
assign addr[6370]= 1380375881;
assign addr[6371]= 1438083551;
assign addr[6372]= 1493966902;
assign addr[6373]= 1547955041;
assign addr[6374]= 1599979481;
assign addr[6375]= 1649974225;
assign addr[6376]= 1697875851;
assign addr[6377]= 1743623590;
assign addr[6378]= 1787159411;
assign addr[6379]= 1828428082;
assign addr[6380]= 1867377253;
assign addr[6381]= 1903957513;
assign addr[6382]= 1938122457;
assign addr[6383]= 1969828744;
assign addr[6384]= 1999036154;
assign addr[6385]= 2025707632;
assign addr[6386]= 2049809346;
assign addr[6387]= 2071310720;
assign addr[6388]= 2090184478;
assign addr[6389]= 2106406677;
assign addr[6390]= 2119956737;
assign addr[6391]= 2130817471;
assign addr[6392]= 2138975100;
assign addr[6393]= 2144419275;
assign addr[6394]= 2147143090;
assign addr[6395]= 2147143090;
assign addr[6396]= 2144419275;
assign addr[6397]= 2138975100;
assign addr[6398]= 2130817471;
assign addr[6399]= 2119956737;
assign addr[6400]= 2106406677;
assign addr[6401]= 2090184478;
assign addr[6402]= 2071310720;
assign addr[6403]= 2049809346;
assign addr[6404]= 2025707632;
assign addr[6405]= 1999036154;
assign addr[6406]= 1969828744;
assign addr[6407]= 1938122457;
assign addr[6408]= 1903957513;
assign addr[6409]= 1867377253;
assign addr[6410]= 1828428082;
assign addr[6411]= 1787159411;
assign addr[6412]= 1743623590;
assign addr[6413]= 1697875851;
assign addr[6414]= 1649974225;
assign addr[6415]= 1599979481;
assign addr[6416]= 1547955041;
assign addr[6417]= 1493966902;
assign addr[6418]= 1438083551;
assign addr[6419]= 1380375881;
assign addr[6420]= 1320917099;
assign addr[6421]= 1259782632;
assign addr[6422]= 1197050035;
assign addr[6423]= 1132798888;
assign addr[6424]= 1067110699;
assign addr[6425]= 1000068799;
assign addr[6426]= 931758235;
assign addr[6427]= 862265664;
assign addr[6428]= 791679244;
assign addr[6429]= 720088517;
assign addr[6430]= 647584304;
assign addr[6431]= 574258580;
assign addr[6432]= 500204365;
assign addr[6433]= 425515602;
assign addr[6434]= 350287041;
assign addr[6435]= 274614114;
assign addr[6436]= 198592817;
assign addr[6437]= 122319591;
assign addr[6438]= 45891193;
assign addr[6439]= -30595422;
assign addr[6440]= -107043224;
assign addr[6441]= -183355234;
assign addr[6442]= -259434643;
assign addr[6443]= -335184940;
assign addr[6444]= -410510029;
assign addr[6445]= -485314355;
assign addr[6446]= -559503022;
assign addr[6447]= -632981917;
assign addr[6448]= -705657826;
assign addr[6449]= -777438554;
assign addr[6450]= -848233042;
assign addr[6451]= -917951481;
assign addr[6452]= -986505429;
assign addr[6453]= -1053807919;
assign addr[6454]= -1119773573;
assign addr[6455]= -1184318708;
assign addr[6456]= -1247361445;
assign addr[6457]= -1308821808;
assign addr[6458]= -1368621831;
assign addr[6459]= -1426685652;
assign addr[6460]= -1482939614;
assign addr[6461]= -1537312353;
assign addr[6462]= -1589734894;
assign addr[6463]= -1640140734;
assign addr[6464]= -1688465931;
assign addr[6465]= -1734649179;
assign addr[6466]= -1778631892;
assign addr[6467]= -1820358275;
assign addr[6468]= -1859775393;
assign addr[6469]= -1896833245;
assign addr[6470]= -1931484818;
assign addr[6471]= -1963686155;
assign addr[6472]= -1993396407;
assign addr[6473]= -2020577882;
assign addr[6474]= -2045196100;
assign addr[6475]= -2067219829;
assign addr[6476]= -2086621133;
assign addr[6477]= -2103375398;
assign addr[6478]= -2117461370;
assign addr[6479]= -2128861181;
assign addr[6480]= -2137560369;
assign addr[6481]= -2143547897;
assign addr[6482]= -2146816171;
assign addr[6483]= -2147361045;
assign addr[6484]= -2145181827;
assign addr[6485]= -2140281282;
assign addr[6486]= -2132665626;
assign addr[6487]= -2122344521;
assign addr[6488]= -2109331059;
assign addr[6489]= -2093641749;
assign addr[6490]= -2075296495;
assign addr[6491]= -2054318569;
assign addr[6492]= -2030734582;
assign addr[6493]= -2004574453;
assign addr[6494]= -1975871368;
assign addr[6495]= -1944661739;
assign addr[6496]= -1910985158;
assign addr[6497]= -1874884346;
assign addr[6498]= -1836405100;
assign addr[6499]= -1795596234;
assign addr[6500]= -1752509516;
assign addr[6501]= -1707199606;
assign addr[6502]= -1659723983;
assign addr[6503]= -1610142873;
assign addr[6504]= -1558519173;
assign addr[6505]= -1504918373;
assign addr[6506]= -1449408469;
assign addr[6507]= -1392059879;
assign addr[6508]= -1332945355;
assign addr[6509]= -1272139887;
assign addr[6510]= -1209720613;
assign addr[6511]= -1145766716;
assign addr[6512]= -1080359326;
assign addr[6513]= -1013581418;
assign addr[6514]= -945517704;
assign addr[6515]= -876254528;
assign addr[6516]= -805879757;
assign addr[6517]= -734482665;
assign addr[6518]= -662153826;
assign addr[6519]= -588984994;
assign addr[6520]= -515068990;
assign addr[6521]= -440499581;
assign addr[6522]= -365371365;
assign addr[6523]= -289779648;
assign addr[6524]= -213820322;
assign addr[6525]= -137589750;
assign addr[6526]= -61184634;
assign addr[6527]= 15298099;
assign addr[6528]= 91761426;
assign addr[6529]= 168108346;
assign addr[6530]= 244242007;
assign addr[6531]= 320065829;
assign addr[6532]= 395483624;
assign addr[6533]= 470399716;
assign addr[6534]= 544719071;
assign addr[6535]= 618347408;
assign addr[6536]= 691191324;
assign addr[6537]= 763158411;
assign addr[6538]= 834157373;
assign addr[6539]= 904098143;
assign addr[6540]= 972891995;
assign addr[6541]= 1040451659;
assign addr[6542]= 1106691431;
assign addr[6543]= 1171527280;
assign addr[6544]= 1234876957;
assign addr[6545]= 1296660098;
assign addr[6546]= 1356798326;
assign addr[6547]= 1415215352;
assign addr[6548]= 1471837070;
assign addr[6549]= 1526591649;
assign addr[6550]= 1579409630;
assign addr[6551]= 1630224009;
assign addr[6552]= 1678970324;
assign addr[6553]= 1725586737;
assign addr[6554]= 1770014111;
assign addr[6555]= 1812196087;
assign addr[6556]= 1852079154;
assign addr[6557]= 1889612716;
assign addr[6558]= 1924749160;
assign addr[6559]= 1957443913;
assign addr[6560]= 1987655498;
assign addr[6561]= 2015345591;
assign addr[6562]= 2040479063;
assign addr[6563]= 2063024031;
assign addr[6564]= 2082951896;
assign addr[6565]= 2100237377;
assign addr[6566]= 2114858546;
assign addr[6567]= 2126796855;
assign addr[6568]= 2136037160;
assign addr[6569]= 2142567738;
assign addr[6570]= 2146380306;
assign addr[6571]= 2147470025;
assign addr[6572]= 2145835515;
assign addr[6573]= 2141478848;
assign addr[6574]= 2134405552;
assign addr[6575]= 2124624598;
assign addr[6576]= 2112148396;
assign addr[6577]= 2096992772;
assign addr[6578]= 2079176953;
assign addr[6579]= 2058723538;
assign addr[6580]= 2035658475;
assign addr[6581]= 2010011024;
assign addr[6582]= 1981813720;
assign addr[6583]= 1951102334;
assign addr[6584]= 1917915825;
assign addr[6585]= 1882296293;
assign addr[6586]= 1844288924;
assign addr[6587]= 1803941934;
assign addr[6588]= 1761306505;
assign addr[6589]= 1716436725;
assign addr[6590]= 1669389513;
assign addr[6591]= 1620224553;
assign addr[6592]= 1569004214;
assign addr[6593]= 1515793473;
assign addr[6594]= 1460659832;
assign addr[6595]= 1403673233;
assign addr[6596]= 1344905966;
assign addr[6597]= 1284432584;
assign addr[6598]= 1222329801;
assign addr[6599]= 1158676398;
assign addr[6600]= 1093553126;
assign addr[6601]= 1027042599;
assign addr[6602]= 959229189;
assign addr[6603]= 890198924;
assign addr[6604]= 820039373;
assign addr[6605]= 748839539;
assign addr[6606]= 676689746;
assign addr[6607]= 603681519;
assign addr[6608]= 529907477;
assign addr[6609]= 455461206;
assign addr[6610]= 380437148;
assign addr[6611]= 304930476;
assign addr[6612]= 229036977;
assign addr[6613]= 152852926;
assign addr[6614]= 76474970;
assign addr[6615]= 0;
assign addr[6616]= -76474970;
assign addr[6617]= -152852926;
assign addr[6618]= -229036977;
assign addr[6619]= -304930476;
assign addr[6620]= -380437148;
assign addr[6621]= -455461206;
assign addr[6622]= -529907477;
assign addr[6623]= -603681519;
assign addr[6624]= -676689746;
assign addr[6625]= -748839539;
assign addr[6626]= -820039373;
assign addr[6627]= -890198924;
assign addr[6628]= -959229189;
assign addr[6629]= -1027042599;
assign addr[6630]= -1093553126;
assign addr[6631]= -1158676398;
assign addr[6632]= -1222329801;
assign addr[6633]= -1284432584;
assign addr[6634]= -1344905966;
assign addr[6635]= -1403673233;
assign addr[6636]= -1460659832;
assign addr[6637]= -1515793473;
assign addr[6638]= -1569004214;
assign addr[6639]= -1620224553;
assign addr[6640]= -1669389513;
assign addr[6641]= -1716436725;
assign addr[6642]= -1761306505;
assign addr[6643]= -1803941934;
assign addr[6644]= -1844288924;
assign addr[6645]= -1882296293;
assign addr[6646]= -1917915825;
assign addr[6647]= -1951102334;
assign addr[6648]= -1981813720;
assign addr[6649]= -2010011024;
assign addr[6650]= -2035658475;
assign addr[6651]= -2058723538;
assign addr[6652]= -2079176953;
assign addr[6653]= -2096992772;
assign addr[6654]= -2112148396;
assign addr[6655]= -2124624598;
assign addr[6656]= -2134405552;
assign addr[6657]= -2141478848;
assign addr[6658]= -2145835515;
assign addr[6659]= -2147470025;
assign addr[6660]= -2146380306;
assign addr[6661]= -2142567738;
assign addr[6662]= -2136037160;
assign addr[6663]= -2126796855;
assign addr[6664]= -2114858546;
assign addr[6665]= -2100237377;
assign addr[6666]= -2082951896;
assign addr[6667]= -2063024031;
assign addr[6668]= -2040479063;
assign addr[6669]= -2015345591;
assign addr[6670]= -1987655498;
assign addr[6671]= -1957443913;
assign addr[6672]= -1924749160;
assign addr[6673]= -1889612716;
assign addr[6674]= -1852079154;
assign addr[6675]= -1812196087;
assign addr[6676]= -1770014111;
assign addr[6677]= -1725586737;
assign addr[6678]= -1678970324;
assign addr[6679]= -1630224009;
assign addr[6680]= -1579409630;
assign addr[6681]= -1526591649;
assign addr[6682]= -1471837070;
assign addr[6683]= -1415215352;
assign addr[6684]= -1356798326;
assign addr[6685]= -1296660098;
assign addr[6686]= -1234876957;
assign addr[6687]= -1171527280;
assign addr[6688]= -1106691431;
assign addr[6689]= -1040451659;
assign addr[6690]= -972891995;
assign addr[6691]= -904098143;
assign addr[6692]= -834157373;
assign addr[6693]= -763158411;
assign addr[6694]= -691191324;
assign addr[6695]= -618347408;
assign addr[6696]= -544719071;
assign addr[6697]= -470399716;
assign addr[6698]= -395483624;
assign addr[6699]= -320065829;
assign addr[6700]= -244242007;
assign addr[6701]= -168108346;
assign addr[6702]= -91761426;
assign addr[6703]= -15298099;
assign addr[6704]= 61184634;
assign addr[6705]= 137589750;
assign addr[6706]= 213820322;
assign addr[6707]= 289779648;
assign addr[6708]= 365371365;
assign addr[6709]= 440499581;
assign addr[6710]= 515068990;
assign addr[6711]= 588984994;
assign addr[6712]= 662153826;
assign addr[6713]= 734482665;
assign addr[6714]= 805879757;
assign addr[6715]= 876254528;
assign addr[6716]= 945517704;
assign addr[6717]= 1013581418;
assign addr[6718]= 1080359326;
assign addr[6719]= 1145766716;
assign addr[6720]= 1209720613;
assign addr[6721]= 1272139887;
assign addr[6722]= 1332945355;
assign addr[6723]= 1392059879;
assign addr[6724]= 1449408469;
assign addr[6725]= 1504918373;
assign addr[6726]= 1558519173;
assign addr[6727]= 1610142873;
assign addr[6728]= 1659723983;
assign addr[6729]= 1707199606;
assign addr[6730]= 1752509516;
assign addr[6731]= 1795596234;
assign addr[6732]= 1836405100;
assign addr[6733]= 1874884346;
assign addr[6734]= 1910985158;
assign addr[6735]= 1944661739;
assign addr[6736]= 1975871368;
assign addr[6737]= 2004574453;
assign addr[6738]= 2030734582;
assign addr[6739]= 2054318569;
assign addr[6740]= 2075296495;
assign addr[6741]= 2093641749;
assign addr[6742]= 2109331059;
assign addr[6743]= 2122344521;
assign addr[6744]= 2132665626;
assign addr[6745]= 2140281282;
assign addr[6746]= 2145181827;
assign addr[6747]= 2147361045;
assign addr[6748]= 2146816171;
assign addr[6749]= 2143547897;
assign addr[6750]= 2137560369;
assign addr[6751]= 2128861181;
assign addr[6752]= 2117461370;
assign addr[6753]= 2103375398;
assign addr[6754]= 2086621133;
assign addr[6755]= 2067219829;
assign addr[6756]= 2045196100;
assign addr[6757]= 2020577882;
assign addr[6758]= 1993396407;
assign addr[6759]= 1963686155;
assign addr[6760]= 1931484818;
assign addr[6761]= 1896833245;
assign addr[6762]= 1859775393;
assign addr[6763]= 1820358275;
assign addr[6764]= 1778631892;
assign addr[6765]= 1734649179;
assign addr[6766]= 1688465931;
assign addr[6767]= 1640140734;
assign addr[6768]= 1589734894;
assign addr[6769]= 1537312353;
assign addr[6770]= 1482939614;
assign addr[6771]= 1426685652;
assign addr[6772]= 1368621831;
assign addr[6773]= 1308821808;
assign addr[6774]= 1247361445;
assign addr[6775]= 1184318708;
assign addr[6776]= 1119773573;
assign addr[6777]= 1053807919;
assign addr[6778]= 986505429;
assign addr[6779]= 917951481;
assign addr[6780]= 848233042;
assign addr[6781]= 777438554;
assign addr[6782]= 705657826;
assign addr[6783]= 632981917;
assign addr[6784]= 559503022;
assign addr[6785]= 485314355;
assign addr[6786]= 410510029;
assign addr[6787]= 335184940;
assign addr[6788]= 259434643;
assign addr[6789]= 183355234;
assign addr[6790]= 107043224;
assign addr[6791]= 30595422;
assign addr[6792]= -45891193;
assign addr[6793]= -122319591;
assign addr[6794]= -198592817;
assign addr[6795]= -274614114;
assign addr[6796]= -350287041;
assign addr[6797]= -425515602;
assign addr[6798]= -500204365;
assign addr[6799]= -574258580;
assign addr[6800]= -647584304;
assign addr[6801]= -720088517;
assign addr[6802]= -791679244;
assign addr[6803]= -862265664;
assign addr[6804]= -931758235;
assign addr[6805]= -1000068799;
assign addr[6806]= -1067110699;
assign addr[6807]= -1132798888;
assign addr[6808]= -1197050035;
assign addr[6809]= -1259782632;
assign addr[6810]= -1320917099;
assign addr[6811]= -1380375881;
assign addr[6812]= -1438083551;
assign addr[6813]= -1493966902;
assign addr[6814]= -1547955041;
assign addr[6815]= -1599979481;
assign addr[6816]= -1649974225;
assign addr[6817]= -1697875851;
assign addr[6818]= -1743623590;
assign addr[6819]= -1787159411;
assign addr[6820]= -1828428082;
assign addr[6821]= -1867377253;
assign addr[6822]= -1903957513;
assign addr[6823]= -1938122457;
assign addr[6824]= -1969828744;
assign addr[6825]= -1999036154;
assign addr[6826]= -2025707632;
assign addr[6827]= -2049809346;
assign addr[6828]= -2071310720;
assign addr[6829]= -2090184478;
assign addr[6830]= -2106406677;
assign addr[6831]= -2119956737;
assign addr[6832]= -2130817471;
assign addr[6833]= -2138975100;
assign addr[6834]= -2144419275;
assign addr[6835]= -2147143090;
assign addr[6836]= -2147143090;
assign addr[6837]= -2144419275;
assign addr[6838]= -2138975100;
assign addr[6839]= -2130817471;
assign addr[6840]= -2119956737;
assign addr[6841]= -2106406677;
assign addr[6842]= -2090184478;
assign addr[6843]= -2071310720;
assign addr[6844]= -2049809346;
assign addr[6845]= -2025707632;
assign addr[6846]= -1999036154;
assign addr[6847]= -1969828744;
assign addr[6848]= -1938122457;
assign addr[6849]= -1903957513;
assign addr[6850]= -1867377253;
assign addr[6851]= -1828428082;
assign addr[6852]= -1787159411;
assign addr[6853]= -1743623590;
assign addr[6854]= -1697875851;
assign addr[6855]= -1649974225;
assign addr[6856]= -1599979481;
assign addr[6857]= -1547955041;
assign addr[6858]= -1493966902;
assign addr[6859]= -1438083551;
assign addr[6860]= -1380375881;
assign addr[6861]= -1320917099;
assign addr[6862]= -1259782632;
assign addr[6863]= -1197050035;
assign addr[6864]= -1132798888;
assign addr[6865]= -1067110699;
assign addr[6866]= -1000068799;
assign addr[6867]= -931758235;
assign addr[6868]= -862265664;
assign addr[6869]= -791679244;
assign addr[6870]= -720088517;
assign addr[6871]= -647584304;
assign addr[6872]= -574258580;
assign addr[6873]= -500204365;
assign addr[6874]= -425515602;
assign addr[6875]= -350287041;
assign addr[6876]= -274614114;
assign addr[6877]= -198592817;
assign addr[6878]= -122319591;
assign addr[6879]= -45891193;
assign addr[6880]= 30595422;
assign addr[6881]= 107043224;
assign addr[6882]= 183355234;
assign addr[6883]= 259434643;
assign addr[6884]= 335184940;
assign addr[6885]= 410510029;
assign addr[6886]= 485314355;
assign addr[6887]= 559503022;
assign addr[6888]= 632981917;
assign addr[6889]= 705657826;
assign addr[6890]= 777438554;
assign addr[6891]= 848233042;
assign addr[6892]= 917951481;
assign addr[6893]= 986505429;
assign addr[6894]= 1053807919;
assign addr[6895]= 1119773573;
assign addr[6896]= 1184318708;
assign addr[6897]= 1247361445;
assign addr[6898]= 1308821808;
assign addr[6899]= 1368621831;
assign addr[6900]= 1426685652;
assign addr[6901]= 1482939614;
assign addr[6902]= 1537312353;
assign addr[6903]= 1589734894;
assign addr[6904]= 1640140734;
assign addr[6905]= 1688465931;
assign addr[6906]= 1734649179;
assign addr[6907]= 1778631892;
assign addr[6908]= 1820358275;
assign addr[6909]= 1859775393;
assign addr[6910]= 1896833245;
assign addr[6911]= 1931484818;
assign addr[6912]= 1963686155;
assign addr[6913]= 1993396407;
assign addr[6914]= 2020577882;
assign addr[6915]= 2045196100;
assign addr[6916]= 2067219829;
assign addr[6917]= 2086621133;
assign addr[6918]= 2103375398;
assign addr[6919]= 2117461370;
assign addr[6920]= 2128861181;
assign addr[6921]= 2137560369;
assign addr[6922]= 2143547897;
assign addr[6923]= 2146816171;
assign addr[6924]= 2147361045;
assign addr[6925]= 2145181827;
assign addr[6926]= 2140281282;
assign addr[6927]= 2132665626;
assign addr[6928]= 2122344521;
assign addr[6929]= 2109331059;
assign addr[6930]= 2093641749;
assign addr[6931]= 2075296495;
assign addr[6932]= 2054318569;
assign addr[6933]= 2030734582;
assign addr[6934]= 2004574453;
assign addr[6935]= 1975871368;
assign addr[6936]= 1944661739;
assign addr[6937]= 1910985158;
assign addr[6938]= 1874884346;
assign addr[6939]= 1836405100;
assign addr[6940]= 1795596234;
assign addr[6941]= 1752509516;
assign addr[6942]= 1707199606;
assign addr[6943]= 1659723983;
assign addr[6944]= 1610142873;
assign addr[6945]= 1558519173;
assign addr[6946]= 1504918373;
assign addr[6947]= 1449408469;
assign addr[6948]= 1392059879;
assign addr[6949]= 1332945355;
assign addr[6950]= 1272139887;
assign addr[6951]= 1209720613;
assign addr[6952]= 1145766716;
assign addr[6953]= 1080359326;
assign addr[6954]= 1013581418;
assign addr[6955]= 945517704;
assign addr[6956]= 876254528;
assign addr[6957]= 805879757;
assign addr[6958]= 734482665;
assign addr[6959]= 662153826;
assign addr[6960]= 588984994;
assign addr[6961]= 515068990;
assign addr[6962]= 440499581;
assign addr[6963]= 365371365;
assign addr[6964]= 289779648;
assign addr[6965]= 213820322;
assign addr[6966]= 137589750;
assign addr[6967]= 61184634;
assign addr[6968]= -15298099;
assign addr[6969]= -91761426;
assign addr[6970]= -168108346;
assign addr[6971]= -244242007;
assign addr[6972]= -320065829;
assign addr[6973]= -395483624;
assign addr[6974]= -470399716;
assign addr[6975]= -544719071;
assign addr[6976]= -618347408;
assign addr[6977]= -691191324;
assign addr[6978]= -763158411;
assign addr[6979]= -834157373;
assign addr[6980]= -904098143;
assign addr[6981]= -972891995;
assign addr[6982]= -1040451659;
assign addr[6983]= -1106691431;
assign addr[6984]= -1171527280;
assign addr[6985]= -1234876957;
assign addr[6986]= -1296660098;
assign addr[6987]= -1356798326;
assign addr[6988]= -1415215352;
assign addr[6989]= -1471837070;
assign addr[6990]= -1526591649;
assign addr[6991]= -1579409630;
assign addr[6992]= -1630224009;
assign addr[6993]= -1678970324;
assign addr[6994]= -1725586737;
assign addr[6995]= -1770014111;
assign addr[6996]= -1812196087;
assign addr[6997]= -1852079154;
assign addr[6998]= -1889612716;
assign addr[6999]= -1924749160;
assign addr[7000]= -1957443913;
assign addr[7001]= -1987655498;
assign addr[7002]= -2015345591;
assign addr[7003]= -2040479063;
assign addr[7004]= -2063024031;
assign addr[7005]= -2082951896;
assign addr[7006]= -2100237377;
assign addr[7007]= -2114858546;
assign addr[7008]= -2126796855;
assign addr[7009]= -2136037160;
assign addr[7010]= -2142567738;
assign addr[7011]= -2146380306;
assign addr[7012]= -2147470025;
assign addr[7013]= -2145835515;
assign addr[7014]= -2141478848;
assign addr[7015]= -2134405552;
assign addr[7016]= -2124624598;
assign addr[7017]= -2112148396;
assign addr[7018]= -2096992772;
assign addr[7019]= -2079176953;
assign addr[7020]= -2058723538;
assign addr[7021]= -2035658475;
assign addr[7022]= -2010011024;
assign addr[7023]= -1981813720;
assign addr[7024]= -1951102334;
assign addr[7025]= -1917915825;
assign addr[7026]= -1882296293;
assign addr[7027]= -1844288924;
assign addr[7028]= -1803941934;
assign addr[7029]= -1761306505;
assign addr[7030]= -1716436725;
assign addr[7031]= -1669389513;
assign addr[7032]= -1620224553;
assign addr[7033]= -1569004214;
assign addr[7034]= -1515793473;
assign addr[7035]= -1460659832;
assign addr[7036]= -1403673233;
assign addr[7037]= -1344905966;
assign addr[7038]= -1284432584;
assign addr[7039]= -1222329801;
assign addr[7040]= -1158676398;
assign addr[7041]= -1093553126;
assign addr[7042]= -1027042599;
assign addr[7043]= -959229189;
assign addr[7044]= -890198924;
assign addr[7045]= -820039373;
assign addr[7046]= -748839539;
assign addr[7047]= -676689746;
assign addr[7048]= -603681519;
assign addr[7049]= -529907477;
assign addr[7050]= -455461206;
assign addr[7051]= -380437148;
assign addr[7052]= -304930476;
assign addr[7053]= -229036977;
assign addr[7054]= -152852926;
assign addr[7055]= -76474970;
assign addr[7056]= 0;
assign addr[7057]= 76474970;
assign addr[7058]= 152852926;
assign addr[7059]= 229036977;
assign addr[7060]= 304930476;
assign addr[7061]= 380437148;
assign addr[7062]= 455461206;
assign addr[7063]= 529907477;
assign addr[7064]= 603681519;
assign addr[7065]= 676689746;
assign addr[7066]= 748839539;
assign addr[7067]= 820039373;
assign addr[7068]= 890198924;
assign addr[7069]= 959229189;
assign addr[7070]= 1027042599;
assign addr[7071]= 1093553126;
assign addr[7072]= 1158676398;
assign addr[7073]= 1222329801;
assign addr[7074]= 1284432584;
assign addr[7075]= 1344905966;
assign addr[7076]= 1403673233;
assign addr[7077]= 1460659832;
assign addr[7078]= 1515793473;
assign addr[7079]= 1569004214;
assign addr[7080]= 1620224553;
assign addr[7081]= 1669389513;
assign addr[7082]= 1716436725;
assign addr[7083]= 1761306505;
assign addr[7084]= 1803941934;
assign addr[7085]= 1844288924;
assign addr[7086]= 1882296293;
assign addr[7087]= 1917915825;
assign addr[7088]= 1951102334;
assign addr[7089]= 1981813720;
assign addr[7090]= 2010011024;
assign addr[7091]= 2035658475;
assign addr[7092]= 2058723538;
assign addr[7093]= 2079176953;
assign addr[7094]= 2096992772;
assign addr[7095]= 2112148396;
assign addr[7096]= 2124624598;
assign addr[7097]= 2134405552;
assign addr[7098]= 2141478848;
assign addr[7099]= 2145835515;
assign addr[7100]= 2147470025;
assign addr[7101]= 2146380306;
assign addr[7102]= 2142567738;
assign addr[7103]= 2136037160;
assign addr[7104]= 2126796855;
assign addr[7105]= 2114858546;
assign addr[7106]= 2100237377;
assign addr[7107]= 2082951896;
assign addr[7108]= 2063024031;
assign addr[7109]= 2040479063;
assign addr[7110]= 2015345591;
assign addr[7111]= 1987655498;
assign addr[7112]= 1957443913;
assign addr[7113]= 1924749160;
assign addr[7114]= 1889612716;
assign addr[7115]= 1852079154;
assign addr[7116]= 1812196087;
assign addr[7117]= 1770014111;
assign addr[7118]= 1725586737;
assign addr[7119]= 1678970324;
assign addr[7120]= 1630224009;
assign addr[7121]= 1579409630;
assign addr[7122]= 1526591649;
assign addr[7123]= 1471837070;
assign addr[7124]= 1415215352;
assign addr[7125]= 1356798326;
assign addr[7126]= 1296660098;
assign addr[7127]= 1234876957;
assign addr[7128]= 1171527280;
assign addr[7129]= 1106691431;
assign addr[7130]= 1040451659;
assign addr[7131]= 972891995;
assign addr[7132]= 904098143;
assign addr[7133]= 834157373;
assign addr[7134]= 763158411;
assign addr[7135]= 691191324;
assign addr[7136]= 618347408;
assign addr[7137]= 544719071;
assign addr[7138]= 470399716;
assign addr[7139]= 395483624;
assign addr[7140]= 320065829;
assign addr[7141]= 244242007;
assign addr[7142]= 168108346;
assign addr[7143]= 91761426;
assign addr[7144]= 15298099;
assign addr[7145]= -61184634;
assign addr[7146]= -137589750;
assign addr[7147]= -213820322;
assign addr[7148]= -289779648;
assign addr[7149]= -365371365;
assign addr[7150]= -440499581;
assign addr[7151]= -515068990;
assign addr[7152]= -588984994;
assign addr[7153]= -662153826;
assign addr[7154]= -734482665;
assign addr[7155]= -805879757;
assign addr[7156]= -876254528;
assign addr[7157]= -945517704;
assign addr[7158]= -1013581418;
assign addr[7159]= -1080359326;
assign addr[7160]= -1145766716;
assign addr[7161]= -1209720613;
assign addr[7162]= -1272139887;
assign addr[7163]= -1332945355;
assign addr[7164]= -1392059879;
assign addr[7165]= -1449408469;
assign addr[7166]= -1504918373;
assign addr[7167]= -1558519173;
assign addr[7168]= -1610142873;
assign addr[7169]= -1659723983;
assign addr[7170]= -1707199606;
assign addr[7171]= -1752509516;
assign addr[7172]= -1795596234;
assign addr[7173]= -1836405100;
assign addr[7174]= -1874884346;
assign addr[7175]= -1910985158;
assign addr[7176]= -1944661739;
assign addr[7177]= -1975871368;
assign addr[7178]= -2004574453;
assign addr[7179]= -2030734582;
assign addr[7180]= -2054318569;
assign addr[7181]= -2075296495;
assign addr[7182]= -2093641749;
assign addr[7183]= -2109331059;
assign addr[7184]= -2122344521;
assign addr[7185]= -2132665626;
assign addr[7186]= -2140281282;
assign addr[7187]= -2145181827;
assign addr[7188]= -2147361045;
assign addr[7189]= -2146816171;
assign addr[7190]= -2143547897;
assign addr[7191]= -2137560369;
assign addr[7192]= -2128861181;
assign addr[7193]= -2117461370;
assign addr[7194]= -2103375398;
assign addr[7195]= -2086621133;
assign addr[7196]= -2067219829;
assign addr[7197]= -2045196100;
assign addr[7198]= -2020577882;
assign addr[7199]= -1993396407;
assign addr[7200]= -1963686155;
assign addr[7201]= -1931484818;
assign addr[7202]= -1896833245;
assign addr[7203]= -1859775393;
assign addr[7204]= -1820358275;
assign addr[7205]= -1778631892;
assign addr[7206]= -1734649179;
assign addr[7207]= -1688465931;
assign addr[7208]= -1640140734;
assign addr[7209]= -1589734894;
assign addr[7210]= -1537312353;
assign addr[7211]= -1482939614;
assign addr[7212]= -1426685652;
assign addr[7213]= -1368621831;
assign addr[7214]= -1308821808;
assign addr[7215]= -1247361445;
assign addr[7216]= -1184318708;
assign addr[7217]= -1119773573;
assign addr[7218]= -1053807919;
assign addr[7219]= -986505429;
assign addr[7220]= -917951481;
assign addr[7221]= -848233042;
assign addr[7222]= -777438554;
assign addr[7223]= -705657826;
assign addr[7224]= -632981917;
assign addr[7225]= -559503022;
assign addr[7226]= -485314355;
assign addr[7227]= -410510029;
assign addr[7228]= -335184940;
assign addr[7229]= -259434643;
assign addr[7230]= -183355234;
assign addr[7231]= -107043224;
assign addr[7232]= -30595422;
assign addr[7233]= 45891193;
assign addr[7234]= 122319591;
assign addr[7235]= 198592817;
assign addr[7236]= 274614114;
assign addr[7237]= 350287041;
assign addr[7238]= 425515602;
assign addr[7239]= 500204365;
assign addr[7240]= 574258580;
assign addr[7241]= 647584304;
assign addr[7242]= 720088517;
assign addr[7243]= 791679244;
assign addr[7244]= 862265664;
assign addr[7245]= 931758235;
assign addr[7246]= 1000068799;
assign addr[7247]= 1067110699;
assign addr[7248]= 1132798888;
assign addr[7249]= 1197050035;
assign addr[7250]= 1259782632;
assign addr[7251]= 1320917099;
assign addr[7252]= 1380375881;
assign addr[7253]= 1438083551;
assign addr[7254]= 1493966902;
assign addr[7255]= 1547955041;
assign addr[7256]= 1599979481;
assign addr[7257]= 1649974225;
assign addr[7258]= 1697875851;
assign addr[7259]= 1743623590;
assign addr[7260]= 1787159411;
assign addr[7261]= 1828428082;
assign addr[7262]= 1867377253;
assign addr[7263]= 1903957513;
assign addr[7264]= 1938122457;
assign addr[7265]= 1969828744;
assign addr[7266]= 1999036154;
assign addr[7267]= 2025707632;
assign addr[7268]= 2049809346;
assign addr[7269]= 2071310720;
assign addr[7270]= 2090184478;
assign addr[7271]= 2106406677;
assign addr[7272]= 2119956737;
assign addr[7273]= 2130817471;
assign addr[7274]= 2138975100;
assign addr[7275]= 2144419275;
assign addr[7276]= 2147143090;
assign addr[7277]= 2147143090;
assign addr[7278]= 2144419275;
assign addr[7279]= 2138975100;
assign addr[7280]= 2130817471;
assign addr[7281]= 2119956737;
assign addr[7282]= 2106406677;
assign addr[7283]= 2090184478;
assign addr[7284]= 2071310720;
assign addr[7285]= 2049809346;
assign addr[7286]= 2025707632;
assign addr[7287]= 1999036154;
assign addr[7288]= 1969828744;
assign addr[7289]= 1938122457;
assign addr[7290]= 1903957513;
assign addr[7291]= 1867377253;
assign addr[7292]= 1828428082;
assign addr[7293]= 1787159411;
assign addr[7294]= 1743623590;
assign addr[7295]= 1697875851;
assign addr[7296]= 1649974225;
assign addr[7297]= 1599979481;
assign addr[7298]= 1547955041;
assign addr[7299]= 1493966902;
assign addr[7300]= 1438083551;
assign addr[7301]= 1380375881;
assign addr[7302]= 1320917099;
assign addr[7303]= 1259782632;
assign addr[7304]= 1197050035;
assign addr[7305]= 1132798888;
assign addr[7306]= 1067110699;
assign addr[7307]= 1000068799;
assign addr[7308]= 931758235;
assign addr[7309]= 862265664;
assign addr[7310]= 791679244;
assign addr[7311]= 720088517;
assign addr[7312]= 647584304;
assign addr[7313]= 574258580;
assign addr[7314]= 500204365;
assign addr[7315]= 425515602;
assign addr[7316]= 350287041;
assign addr[7317]= 274614114;
assign addr[7318]= 198592817;
assign addr[7319]= 122319591;
assign addr[7320]= 45891193;
assign addr[7321]= -30595422;
assign addr[7322]= -107043224;
assign addr[7323]= -183355234;
assign addr[7324]= -259434643;
assign addr[7325]= -335184940;
assign addr[7326]= -410510029;
assign addr[7327]= -485314355;
assign addr[7328]= -559503022;
assign addr[7329]= -632981917;
assign addr[7330]= -705657826;
assign addr[7331]= -777438554;
assign addr[7332]= -848233042;
assign addr[7333]= -917951481;
assign addr[7334]= -986505429;
assign addr[7335]= -1053807919;
assign addr[7336]= -1119773573;
assign addr[7337]= -1184318708;
assign addr[7338]= -1247361445;
assign addr[7339]= -1308821808;
assign addr[7340]= -1368621831;
assign addr[7341]= -1426685652;
assign addr[7342]= -1482939614;
assign addr[7343]= -1537312353;
assign addr[7344]= -1589734894;
assign addr[7345]= -1640140734;
assign addr[7346]= -1688465931;
assign addr[7347]= -1734649179;
assign addr[7348]= -1778631892;
assign addr[7349]= -1820358275;
assign addr[7350]= -1859775393;
assign addr[7351]= -1896833245;
assign addr[7352]= -1931484818;
assign addr[7353]= -1963686155;
assign addr[7354]= -1993396407;
assign addr[7355]= -2020577882;
assign addr[7356]= -2045196100;
assign addr[7357]= -2067219829;
assign addr[7358]= -2086621133;
assign addr[7359]= -2103375398;
assign addr[7360]= -2117461370;
assign addr[7361]= -2128861181;
assign addr[7362]= -2137560369;
assign addr[7363]= -2143547897;
assign addr[7364]= -2146816171;
assign addr[7365]= -2147361045;
assign addr[7366]= -2145181827;
assign addr[7367]= -2140281282;
assign addr[7368]= -2132665626;
assign addr[7369]= -2122344521;
assign addr[7370]= -2109331059;
assign addr[7371]= -2093641749;
assign addr[7372]= -2075296495;
assign addr[7373]= -2054318569;
assign addr[7374]= -2030734582;
assign addr[7375]= -2004574453;
assign addr[7376]= -1975871368;
assign addr[7377]= -1944661739;
assign addr[7378]= -1910985158;
assign addr[7379]= -1874884346;
assign addr[7380]= -1836405100;
assign addr[7381]= -1795596234;
assign addr[7382]= -1752509516;
assign addr[7383]= -1707199606;
assign addr[7384]= -1659723983;
assign addr[7385]= -1610142873;
assign addr[7386]= -1558519173;
assign addr[7387]= -1504918373;
assign addr[7388]= -1449408469;
assign addr[7389]= -1392059879;
assign addr[7390]= -1332945355;
assign addr[7391]= -1272139887;
assign addr[7392]= -1209720613;
assign addr[7393]= -1145766716;
assign addr[7394]= -1080359326;
assign addr[7395]= -1013581418;
assign addr[7396]= -945517704;
assign addr[7397]= -876254528;
assign addr[7398]= -805879757;
assign addr[7399]= -734482665;
assign addr[7400]= -662153826;
assign addr[7401]= -588984994;
assign addr[7402]= -515068990;
assign addr[7403]= -440499581;
assign addr[7404]= -365371365;
assign addr[7405]= -289779648;
assign addr[7406]= -213820322;
assign addr[7407]= -137589750;
assign addr[7408]= -61184634;
assign addr[7409]= 15298099;
assign addr[7410]= 91761426;
assign addr[7411]= 168108346;
assign addr[7412]= 244242007;
assign addr[7413]= 320065829;
assign addr[7414]= 395483624;
assign addr[7415]= 470399716;
assign addr[7416]= 544719071;
assign addr[7417]= 618347408;
assign addr[7418]= 691191324;
assign addr[7419]= 763158411;
assign addr[7420]= 834157373;
assign addr[7421]= 904098143;
assign addr[7422]= 972891995;
assign addr[7423]= 1040451659;
assign addr[7424]= 1106691431;
assign addr[7425]= 1171527280;
assign addr[7426]= 1234876957;
assign addr[7427]= 1296660098;
assign addr[7428]= 1356798326;
assign addr[7429]= 1415215352;
assign addr[7430]= 1471837070;
assign addr[7431]= 1526591649;
assign addr[7432]= 1579409630;
assign addr[7433]= 1630224009;
assign addr[7434]= 1678970324;
assign addr[7435]= 1725586737;
assign addr[7436]= 1770014111;
assign addr[7437]= 1812196087;
assign addr[7438]= 1852079154;
assign addr[7439]= 1889612716;
assign addr[7440]= 1924749160;
assign addr[7441]= 1957443913;
assign addr[7442]= 1987655498;
assign addr[7443]= 2015345591;
assign addr[7444]= 2040479063;
assign addr[7445]= 2063024031;
assign addr[7446]= 2082951896;
assign addr[7447]= 2100237377;
assign addr[7448]= 2114858546;
assign addr[7449]= 2126796855;
assign addr[7450]= 2136037160;
assign addr[7451]= 2142567738;
assign addr[7452]= 2146380306;
assign addr[7453]= 2147470025;
assign addr[7454]= 2145835515;
assign addr[7455]= 2141478848;
assign addr[7456]= 2134405552;
assign addr[7457]= 2124624598;
assign addr[7458]= 2112148396;
assign addr[7459]= 2096992772;
assign addr[7460]= 2079176953;
assign addr[7461]= 2058723538;
assign addr[7462]= 2035658475;
assign addr[7463]= 2010011024;
assign addr[7464]= 1981813720;
assign addr[7465]= 1951102334;
assign addr[7466]= 1917915825;
assign addr[7467]= 1882296293;
assign addr[7468]= 1844288924;
assign addr[7469]= 1803941934;
assign addr[7470]= 1761306505;
assign addr[7471]= 1716436725;
assign addr[7472]= 1669389513;
assign addr[7473]= 1620224553;
assign addr[7474]= 1569004214;
assign addr[7475]= 1515793473;
assign addr[7476]= 1460659832;
assign addr[7477]= 1403673233;
assign addr[7478]= 1344905966;
assign addr[7479]= 1284432584;
assign addr[7480]= 1222329801;
assign addr[7481]= 1158676398;
assign addr[7482]= 1093553126;
assign addr[7483]= 1027042599;
assign addr[7484]= 959229189;
assign addr[7485]= 890198924;
assign addr[7486]= 820039373;
assign addr[7487]= 748839539;
assign addr[7488]= 676689746;
assign addr[7489]= 603681519;
assign addr[7490]= 529907477;
assign addr[7491]= 455461206;
assign addr[7492]= 380437148;
assign addr[7493]= 304930476;
assign addr[7494]= 229036977;
assign addr[7495]= 152852926;
assign addr[7496]= 76474970;
assign addr[7497]= 0;
assign addr[7498]= -76474970;
assign addr[7499]= -152852926;
assign addr[7500]= -229036977;
assign addr[7501]= -304930476;
assign addr[7502]= -380437148;
assign addr[7503]= -455461206;
assign addr[7504]= -529907477;
assign addr[7505]= -603681519;
assign addr[7506]= -676689746;
assign addr[7507]= -748839539;
assign addr[7508]= -820039373;
assign addr[7509]= -890198924;
assign addr[7510]= -959229189;
assign addr[7511]= -1027042599;
assign addr[7512]= -1093553126;
assign addr[7513]= -1158676398;
assign addr[7514]= -1222329801;
assign addr[7515]= -1284432584;
assign addr[7516]= -1344905966;
assign addr[7517]= -1403673233;
assign addr[7518]= -1460659832;
assign addr[7519]= -1515793473;
assign addr[7520]= -1569004214;
assign addr[7521]= -1620224553;
assign addr[7522]= -1669389513;
assign addr[7523]= -1716436725;
assign addr[7524]= -1761306505;
assign addr[7525]= -1803941934;
assign addr[7526]= -1844288924;
assign addr[7527]= -1882296293;
assign addr[7528]= -1917915825;
assign addr[7529]= -1951102334;
assign addr[7530]= -1981813720;
assign addr[7531]= -2010011024;
assign addr[7532]= -2035658475;
assign addr[7533]= -2058723538;
assign addr[7534]= -2079176953;
assign addr[7535]= -2096992772;
assign addr[7536]= -2112148396;
assign addr[7537]= -2124624598;
assign addr[7538]= -2134405552;
assign addr[7539]= -2141478848;
assign addr[7540]= -2145835515;
assign addr[7541]= -2147470025;
assign addr[7542]= -2146380306;
assign addr[7543]= -2142567738;
assign addr[7544]= -2136037160;
assign addr[7545]= -2126796855;
assign addr[7546]= -2114858546;
assign addr[7547]= -2100237377;
assign addr[7548]= -2082951896;
assign addr[7549]= -2063024031;
assign addr[7550]= -2040479063;
assign addr[7551]= -2015345591;
assign addr[7552]= -1987655498;
assign addr[7553]= -1957443913;
assign addr[7554]= -1924749160;
assign addr[7555]= -1889612716;
assign addr[7556]= -1852079154;
assign addr[7557]= -1812196087;
assign addr[7558]= -1770014111;
assign addr[7559]= -1725586737;
assign addr[7560]= -1678970324;
assign addr[7561]= -1630224009;
assign addr[7562]= -1579409630;
assign addr[7563]= -1526591649;
assign addr[7564]= -1471837070;
assign addr[7565]= -1415215352;
assign addr[7566]= -1356798326;
assign addr[7567]= -1296660098;
assign addr[7568]= -1234876957;
assign addr[7569]= -1171527280;
assign addr[7570]= -1106691431;
assign addr[7571]= -1040451659;
assign addr[7572]= -972891995;
assign addr[7573]= -904098143;
assign addr[7574]= -834157373;
assign addr[7575]= -763158411;
assign addr[7576]= -691191324;
assign addr[7577]= -618347408;
assign addr[7578]= -544719071;
assign addr[7579]= -470399716;
assign addr[7580]= -395483624;
assign addr[7581]= -320065829;
assign addr[7582]= -244242007;
assign addr[7583]= -168108346;
assign addr[7584]= -91761426;
assign addr[7585]= -15298099;
assign addr[7586]= 61184634;
assign addr[7587]= 137589750;
assign addr[7588]= 213820322;
assign addr[7589]= 289779648;
assign addr[7590]= 365371365;
assign addr[7591]= 440499581;
assign addr[7592]= 515068990;
assign addr[7593]= 588984994;
assign addr[7594]= 662153826;
assign addr[7595]= 734482665;
assign addr[7596]= 805879757;
assign addr[7597]= 876254528;
assign addr[7598]= 945517704;
assign addr[7599]= 1013581418;
assign addr[7600]= 1080359326;
assign addr[7601]= 1145766716;
assign addr[7602]= 1209720613;
assign addr[7603]= 1272139887;
assign addr[7604]= 1332945355;
assign addr[7605]= 1392059879;
assign addr[7606]= 1449408469;
assign addr[7607]= 1504918373;
assign addr[7608]= 1558519173;
assign addr[7609]= 1610142873;
assign addr[7610]= 1659723983;
assign addr[7611]= 1707199606;
assign addr[7612]= 1752509516;
assign addr[7613]= 1795596234;
assign addr[7614]= 1836405100;
assign addr[7615]= 1874884346;
assign addr[7616]= 1910985158;
assign addr[7617]= 1944661739;
assign addr[7618]= 1975871368;
assign addr[7619]= 2004574453;
assign addr[7620]= 2030734582;
assign addr[7621]= 2054318569;
assign addr[7622]= 2075296495;
assign addr[7623]= 2093641749;
assign addr[7624]= 2109331059;
assign addr[7625]= 2122344521;
assign addr[7626]= 2132665626;
assign addr[7627]= 2140281282;
assign addr[7628]= 2145181827;
assign addr[7629]= 2147361045;
assign addr[7630]= 2146816171;
assign addr[7631]= 2143547897;
assign addr[7632]= 2137560369;
assign addr[7633]= 2128861181;
assign addr[7634]= 2117461370;
assign addr[7635]= 2103375398;
assign addr[7636]= 2086621133;
assign addr[7637]= 2067219829;
assign addr[7638]= 2045196100;
assign addr[7639]= 2020577882;
assign addr[7640]= 1993396407;
assign addr[7641]= 1963686155;
assign addr[7642]= 1931484818;
assign addr[7643]= 1896833245;
assign addr[7644]= 1859775393;
assign addr[7645]= 1820358275;
assign addr[7646]= 1778631892;
assign addr[7647]= 1734649179;
assign addr[7648]= 1688465931;
assign addr[7649]= 1640140734;
assign addr[7650]= 1589734894;
assign addr[7651]= 1537312353;
assign addr[7652]= 1482939614;
assign addr[7653]= 1426685652;
assign addr[7654]= 1368621831;
assign addr[7655]= 1308821808;
assign addr[7656]= 1247361445;
assign addr[7657]= 1184318708;
assign addr[7658]= 1119773573;
assign addr[7659]= 1053807919;
assign addr[7660]= 986505429;
assign addr[7661]= 917951481;
assign addr[7662]= 848233042;
assign addr[7663]= 777438554;
assign addr[7664]= 705657826;
assign addr[7665]= 632981917;
assign addr[7666]= 559503022;
assign addr[7667]= 485314355;
assign addr[7668]= 410510029;
assign addr[7669]= 335184940;
assign addr[7670]= 259434643;
assign addr[7671]= 183355234;
assign addr[7672]= 107043224;
assign addr[7673]= 30595422;
assign addr[7674]= -45891193;
assign addr[7675]= -122319591;
assign addr[7676]= -198592817;
assign addr[7677]= -274614114;
assign addr[7678]= -350287041;
assign addr[7679]= -425515602;
assign addr[7680]= -500204365;
assign addr[7681]= -574258580;
assign addr[7682]= -647584304;
assign addr[7683]= -720088517;
assign addr[7684]= -791679244;
assign addr[7685]= -862265664;
assign addr[7686]= -931758235;
assign addr[7687]= -1000068799;
assign addr[7688]= -1067110699;
assign addr[7689]= -1132798888;
assign addr[7690]= -1197050035;
assign addr[7691]= -1259782632;
assign addr[7692]= -1320917099;
assign addr[7693]= -1380375881;
assign addr[7694]= -1438083551;
assign addr[7695]= -1493966902;
assign addr[7696]= -1547955041;
assign addr[7697]= -1599979481;
assign addr[7698]= -1649974225;
assign addr[7699]= -1697875851;
assign addr[7700]= -1743623590;
assign addr[7701]= -1787159411;
assign addr[7702]= -1828428082;
assign addr[7703]= -1867377253;
assign addr[7704]= -1903957513;
assign addr[7705]= -1938122457;
assign addr[7706]= -1969828744;
assign addr[7707]= -1999036154;
assign addr[7708]= -2025707632;
assign addr[7709]= -2049809346;
assign addr[7710]= -2071310720;
assign addr[7711]= -2090184478;
assign addr[7712]= -2106406677;
assign addr[7713]= -2119956737;
assign addr[7714]= -2130817471;
assign addr[7715]= -2138975100;
assign addr[7716]= -2144419275;
assign addr[7717]= -2147143090;
assign addr[7718]= -2147143090;
assign addr[7719]= -2144419275;
assign addr[7720]= -2138975100;
assign addr[7721]= -2130817471;
assign addr[7722]= -2119956737;
assign addr[7723]= -2106406677;
assign addr[7724]= -2090184478;
assign addr[7725]= -2071310720;
assign addr[7726]= -2049809346;
assign addr[7727]= -2025707632;
assign addr[7728]= -1999036154;
assign addr[7729]= -1969828744;
assign addr[7730]= -1938122457;
assign addr[7731]= -1903957513;
assign addr[7732]= -1867377253;
assign addr[7733]= -1828428082;
assign addr[7734]= -1787159411;
assign addr[7735]= -1743623590;
assign addr[7736]= -1697875851;
assign addr[7737]= -1649974225;
assign addr[7738]= -1599979481;
assign addr[7739]= -1547955041;
assign addr[7740]= -1493966902;
assign addr[7741]= -1438083551;
assign addr[7742]= -1380375881;
assign addr[7743]= -1320917099;
assign addr[7744]= -1259782632;
assign addr[7745]= -1197050035;
assign addr[7746]= -1132798888;
assign addr[7747]= -1067110699;
assign addr[7748]= -1000068799;
assign addr[7749]= -931758235;
assign addr[7750]= -862265664;
assign addr[7751]= -791679244;
assign addr[7752]= -720088517;
assign addr[7753]= -647584304;
assign addr[7754]= -574258580;
assign addr[7755]= -500204365;
assign addr[7756]= -425515602;
assign addr[7757]= -350287041;
assign addr[7758]= -274614114;
assign addr[7759]= -198592817;
assign addr[7760]= -122319591;
assign addr[7761]= -45891193;
assign addr[7762]= 30595422;
assign addr[7763]= 107043224;
assign addr[7764]= 183355234;
assign addr[7765]= 259434643;
assign addr[7766]= 335184940;
assign addr[7767]= 410510029;
assign addr[7768]= 485314355;
assign addr[7769]= 559503022;
assign addr[7770]= 632981917;
assign addr[7771]= 705657826;
assign addr[7772]= 777438554;
assign addr[7773]= 848233042;
assign addr[7774]= 917951481;
assign addr[7775]= 986505429;
assign addr[7776]= 1053807919;
assign addr[7777]= 1119773573;
assign addr[7778]= 1184318708;
assign addr[7779]= 1247361445;
assign addr[7780]= 1308821808;
assign addr[7781]= 1368621831;
assign addr[7782]= 1426685652;
assign addr[7783]= 1482939614;
assign addr[7784]= 1537312353;
assign addr[7785]= 1589734894;
assign addr[7786]= 1640140734;
assign addr[7787]= 1688465931;
assign addr[7788]= 1734649179;
assign addr[7789]= 1778631892;
assign addr[7790]= 1820358275;
assign addr[7791]= 1859775393;
assign addr[7792]= 1896833245;
assign addr[7793]= 1931484818;
assign addr[7794]= 1963686155;
assign addr[7795]= 1993396407;
assign addr[7796]= 2020577882;
assign addr[7797]= 2045196100;
assign addr[7798]= 2067219829;
assign addr[7799]= 2086621133;
assign addr[7800]= 2103375398;
assign addr[7801]= 2117461370;
assign addr[7802]= 2128861181;
assign addr[7803]= 2137560369;
assign addr[7804]= 2143547897;
assign addr[7805]= 2146816171;
assign addr[7806]= 2147361045;
assign addr[7807]= 2145181827;
assign addr[7808]= 2140281282;
assign addr[7809]= 2132665626;
assign addr[7810]= 2122344521;
assign addr[7811]= 2109331059;
assign addr[7812]= 2093641749;
assign addr[7813]= 2075296495;
assign addr[7814]= 2054318569;
assign addr[7815]= 2030734582;
assign addr[7816]= 2004574453;
assign addr[7817]= 1975871368;
assign addr[7818]= 1944661739;
assign addr[7819]= 1910985158;
assign addr[7820]= 1874884346;
assign addr[7821]= 1836405100;
assign addr[7822]= 1795596234;
assign addr[7823]= 1752509516;
assign addr[7824]= 1707199606;
assign addr[7825]= 1659723983;
assign addr[7826]= 1610142873;
assign addr[7827]= 1558519173;
assign addr[7828]= 1504918373;
assign addr[7829]= 1449408469;
assign addr[7830]= 1392059879;
assign addr[7831]= 1332945355;
assign addr[7832]= 1272139887;
assign addr[7833]= 1209720613;
assign addr[7834]= 1145766716;
assign addr[7835]= 1080359326;
assign addr[7836]= 1013581418;
assign addr[7837]= 945517704;
assign addr[7838]= 876254528;
assign addr[7839]= 805879757;
assign addr[7840]= 734482665;
assign addr[7841]= 662153826;
assign addr[7842]= 588984994;
assign addr[7843]= 515068990;
assign addr[7844]= 440499581;
assign addr[7845]= 365371365;
assign addr[7846]= 289779648;
assign addr[7847]= 213820322;
assign addr[7848]= 137589750;
assign addr[7849]= 61184634;
assign addr[7850]= -15298099;
assign addr[7851]= -91761426;
assign addr[7852]= -168108346;
assign addr[7853]= -244242007;
assign addr[7854]= -320065829;
assign addr[7855]= -395483624;
assign addr[7856]= -470399716;
assign addr[7857]= -544719071;
assign addr[7858]= -618347408;
assign addr[7859]= -691191324;
assign addr[7860]= -763158411;
assign addr[7861]= -834157373;
assign addr[7862]= -904098143;
assign addr[7863]= -972891995;
assign addr[7864]= -1040451659;
assign addr[7865]= -1106691431;
assign addr[7866]= -1171527280;
assign addr[7867]= -1234876957;
assign addr[7868]= -1296660098;
assign addr[7869]= -1356798326;
assign addr[7870]= -1415215352;
assign addr[7871]= -1471837070;
assign addr[7872]= -1526591649;
assign addr[7873]= -1579409630;
assign addr[7874]= -1630224009;
assign addr[7875]= -1678970324;
assign addr[7876]= -1725586737;
assign addr[7877]= -1770014111;
assign addr[7878]= -1812196087;
assign addr[7879]= -1852079154;
assign addr[7880]= -1889612716;
assign addr[7881]= -1924749160;
assign addr[7882]= -1957443913;
assign addr[7883]= -1987655498;
assign addr[7884]= -2015345591;
assign addr[7885]= -2040479063;
assign addr[7886]= -2063024031;
assign addr[7887]= -2082951896;
assign addr[7888]= -2100237377;
assign addr[7889]= -2114858546;
assign addr[7890]= -2126796855;
assign addr[7891]= -2136037160;
assign addr[7892]= -2142567738;
assign addr[7893]= -2146380306;
assign addr[7894]= -2147470025;
assign addr[7895]= -2145835515;
assign addr[7896]= -2141478848;
assign addr[7897]= -2134405552;
assign addr[7898]= -2124624598;
assign addr[7899]= -2112148396;
assign addr[7900]= -2096992772;
assign addr[7901]= -2079176953;
assign addr[7902]= -2058723538;
assign addr[7903]= -2035658475;
assign addr[7904]= -2010011024;
assign addr[7905]= -1981813720;
assign addr[7906]= -1951102334;
assign addr[7907]= -1917915825;
assign addr[7908]= -1882296293;
assign addr[7909]= -1844288924;
assign addr[7910]= -1803941934;
assign addr[7911]= -1761306505;
assign addr[7912]= -1716436725;
assign addr[7913]= -1669389513;
assign addr[7914]= -1620224553;
assign addr[7915]= -1569004214;
assign addr[7916]= -1515793473;
assign addr[7917]= -1460659832;
assign addr[7918]= -1403673233;
assign addr[7919]= -1344905966;
assign addr[7920]= -1284432584;
assign addr[7921]= -1222329801;
assign addr[7922]= -1158676398;
assign addr[7923]= -1093553126;
assign addr[7924]= -1027042599;
assign addr[7925]= -959229189;
assign addr[7926]= -890198924;
assign addr[7927]= -820039373;
assign addr[7928]= -748839539;
assign addr[7929]= -676689746;
assign addr[7930]= -603681519;
assign addr[7931]= -529907477;
assign addr[7932]= -455461206;
assign addr[7933]= -380437148;
assign addr[7934]= -304930476;
assign addr[7935]= -229036977;
assign addr[7936]= -152852926;
assign addr[7937]= -76474970;
assign addr[7938]= 0;
assign addr[7939]= 76474970;
assign addr[7940]= 152852926;
assign addr[7941]= 229036977;
assign addr[7942]= 304930476;
assign addr[7943]= 380437148;
assign addr[7944]= 455461206;
assign addr[7945]= 529907477;
assign addr[7946]= 603681519;
assign addr[7947]= 676689746;
assign addr[7948]= 748839539;
assign addr[7949]= 820039373;
assign addr[7950]= 890198924;
assign addr[7951]= 959229189;
assign addr[7952]= 1027042599;
assign addr[7953]= 1093553126;
assign addr[7954]= 1158676398;
assign addr[7955]= 1222329801;
assign addr[7956]= 1284432584;
assign addr[7957]= 1344905966;
assign addr[7958]= 1403673233;
assign addr[7959]= 1460659832;
assign addr[7960]= 1515793473;
assign addr[7961]= 1569004214;
assign addr[7962]= 1620224553;
assign addr[7963]= 1669389513;
assign addr[7964]= 1716436725;
assign addr[7965]= 1761306505;
assign addr[7966]= 1803941934;
assign addr[7967]= 1844288924;
assign addr[7968]= 1882296293;
assign addr[7969]= 1917915825;
assign addr[7970]= 1951102334;
assign addr[7971]= 1981813720;
assign addr[7972]= 2010011024;
assign addr[7973]= 2035658475;
assign addr[7974]= 2058723538;
assign addr[7975]= 2079176953;
assign addr[7976]= 2096992772;
assign addr[7977]= 2112148396;
assign addr[7978]= 2124624598;
assign addr[7979]= 2134405552;
assign addr[7980]= 2141478848;
assign addr[7981]= 2145835515;
assign addr[7982]= 2147470025;
assign addr[7983]= 2146380306;
assign addr[7984]= 2142567738;
assign addr[7985]= 2136037160;
assign addr[7986]= 2126796855;
assign addr[7987]= 2114858546;
assign addr[7988]= 2100237377;
assign addr[7989]= 2082951896;
assign addr[7990]= 2063024031;
assign addr[7991]= 2040479063;
assign addr[7992]= 2015345591;
assign addr[7993]= 1987655498;
assign addr[7994]= 1957443913;
assign addr[7995]= 1924749160;
assign addr[7996]= 1889612716;
assign addr[7997]= 1852079154;
assign addr[7998]= 1812196087;
assign addr[7999]= 1770014111;
assign addr[8000]= 1725586737;
assign addr[8001]= 1678970324;
assign addr[8002]= 1630224009;
assign addr[8003]= 1579409630;
assign addr[8004]= 1526591649;
assign addr[8005]= 1471837070;
assign addr[8006]= 1415215352;
assign addr[8007]= 1356798326;
assign addr[8008]= 1296660098;
assign addr[8009]= 1234876957;
assign addr[8010]= 1171527280;
assign addr[8011]= 1106691431;
assign addr[8012]= 1040451659;
assign addr[8013]= 972891995;
assign addr[8014]= 904098143;
assign addr[8015]= 834157373;
assign addr[8016]= 763158411;
assign addr[8017]= 691191324;
assign addr[8018]= 618347408;
assign addr[8019]= 544719071;
assign addr[8020]= 470399716;
assign addr[8021]= 395483624;
assign addr[8022]= 320065829;
assign addr[8023]= 244242007;
assign addr[8024]= 168108346;
assign addr[8025]= 91761426;
assign addr[8026]= 15298099;
assign addr[8027]= -61184634;
assign addr[8028]= -137589750;
assign addr[8029]= -213820322;
assign addr[8030]= -289779648;
assign addr[8031]= -365371365;
assign addr[8032]= -440499581;
assign addr[8033]= -515068990;
assign addr[8034]= -588984994;
assign addr[8035]= -662153826;
assign addr[8036]= -734482665;
assign addr[8037]= -805879757;
assign addr[8038]= -876254528;
assign addr[8039]= -945517704;
assign addr[8040]= -1013581418;
assign addr[8041]= -1080359326;
assign addr[8042]= -1145766716;
assign addr[8043]= -1209720613;
assign addr[8044]= -1272139887;
assign addr[8045]= -1332945355;
assign addr[8046]= -1392059879;
assign addr[8047]= -1449408469;
assign addr[8048]= -1504918373;
assign addr[8049]= -1558519173;
assign addr[8050]= -1610142873;
assign addr[8051]= -1659723983;
assign addr[8052]= -1707199606;
assign addr[8053]= -1752509516;
assign addr[8054]= -1795596234;
assign addr[8055]= -1836405100;
assign addr[8056]= -1874884346;
assign addr[8057]= -1910985158;
assign addr[8058]= -1944661739;
assign addr[8059]= -1975871368;
assign addr[8060]= -2004574453;
assign addr[8061]= -2030734582;
assign addr[8062]= -2054318569;
assign addr[8063]= -2075296495;
assign addr[8064]= -2093641749;
assign addr[8065]= -2109331059;
assign addr[8066]= -2122344521;
assign addr[8067]= -2132665626;
assign addr[8068]= -2140281282;
assign addr[8069]= -2145181827;
assign addr[8070]= -2147361045;
assign addr[8071]= -2146816171;
assign addr[8072]= -2143547897;
assign addr[8073]= -2137560369;
assign addr[8074]= -2128861181;
assign addr[8075]= -2117461370;
assign addr[8076]= -2103375398;
assign addr[8077]= -2086621133;
assign addr[8078]= -2067219829;
assign addr[8079]= -2045196100;
assign addr[8080]= -2020577882;
assign addr[8081]= -1993396407;
assign addr[8082]= -1963686155;
assign addr[8083]= -1931484818;
assign addr[8084]= -1896833245;
assign addr[8085]= -1859775393;
assign addr[8086]= -1820358275;
assign addr[8087]= -1778631892;
assign addr[8088]= -1734649179;
assign addr[8089]= -1688465931;
assign addr[8090]= -1640140734;
assign addr[8091]= -1589734894;
assign addr[8092]= -1537312353;
assign addr[8093]= -1482939614;
assign addr[8094]= -1426685652;
assign addr[8095]= -1368621831;
assign addr[8096]= -1308821808;
assign addr[8097]= -1247361445;
assign addr[8098]= -1184318708;
assign addr[8099]= -1119773573;
assign addr[8100]= -1053807919;
assign addr[8101]= -986505429;
assign addr[8102]= -917951481;
assign addr[8103]= -848233042;
assign addr[8104]= -777438554;
assign addr[8105]= -705657826;
assign addr[8106]= -632981917;
assign addr[8107]= -559503022;
assign addr[8108]= -485314355;
assign addr[8109]= -410510029;
assign addr[8110]= -335184940;
assign addr[8111]= -259434643;
assign addr[8112]= -183355234;
assign addr[8113]= -107043224;
assign addr[8114]= -30595422;
assign addr[8115]= 45891193;
assign addr[8116]= 122319591;
assign addr[8117]= 198592817;
assign addr[8118]= 274614114;
assign addr[8119]= 350287041;
assign addr[8120]= 425515602;
assign addr[8121]= 500204365;
assign addr[8122]= 574258580;
assign addr[8123]= 647584304;
assign addr[8124]= 720088517;
assign addr[8125]= 791679244;
assign addr[8126]= 862265664;
assign addr[8127]= 931758235;
assign addr[8128]= 1000068799;
assign addr[8129]= 1067110699;
assign addr[8130]= 1132798888;
assign addr[8131]= 1197050035;
assign addr[8132]= 1259782632;
assign addr[8133]= 1320917099;
assign addr[8134]= 1380375881;
assign addr[8135]= 1438083551;
assign addr[8136]= 1493966902;
assign addr[8137]= 1547955041;
assign addr[8138]= 1599979481;
assign addr[8139]= 1649974225;
assign addr[8140]= 1697875851;
assign addr[8141]= 1743623590;
assign addr[8142]= 1787159411;
assign addr[8143]= 1828428082;
assign addr[8144]= 1867377253;
assign addr[8145]= 1903957513;
assign addr[8146]= 1938122457;
assign addr[8147]= 1969828744;
assign addr[8148]= 1999036154;
assign addr[8149]= 2025707632;
assign addr[8150]= 2049809346;
assign addr[8151]= 2071310720;
assign addr[8152]= 2090184478;
assign addr[8153]= 2106406677;
assign addr[8154]= 2119956737;
assign addr[8155]= 2130817471;
assign addr[8156]= 2138975100;
assign addr[8157]= 2144419275;
assign addr[8158]= 2147143090;
assign addr[8159]= 2147143090;
assign addr[8160]= 2144419275;
assign addr[8161]= 2138975100;
assign addr[8162]= 2130817471;
assign addr[8163]= 2119956737;
assign addr[8164]= 2106406677;
assign addr[8165]= 2090184478;
assign addr[8166]= 2071310720;
assign addr[8167]= 2049809346;
assign addr[8168]= 2025707632;
assign addr[8169]= 1999036154;
assign addr[8170]= 1969828744;
assign addr[8171]= 1938122457;
assign addr[8172]= 1903957513;
assign addr[8173]= 1867377253;
assign addr[8174]= 1828428082;
assign addr[8175]= 1787159411;
assign addr[8176]= 1743623590;
assign addr[8177]= 1697875851;
assign addr[8178]= 1649974225;
assign addr[8179]= 1599979481;
assign addr[8180]= 1547955041;
assign addr[8181]= 1493966902;
assign addr[8182]= 1438083551;
assign addr[8183]= 1380375881;
assign addr[8184]= 1320917099;
assign addr[8185]= 1259782632;
assign addr[8186]= 1197050035;
assign addr[8187]= 1132798888;
assign addr[8188]= 1067110699;
assign addr[8189]= 1000068799;
assign addr[8190]= 931758235;
assign addr[8191]= 862265664;
assign addr[8192]= 791679244;
assign addr[8193]= 720088517;
assign addr[8194]= 647584304;
assign addr[8195]= 574258580;
assign addr[8196]= 500204365;
assign addr[8197]= 425515602;
assign addr[8198]= 350287041;
assign addr[8199]= 274614114;
assign addr[8200]= 198592817;
assign addr[8201]= 122319591;
assign addr[8202]= 45891193;
assign addr[8203]= -30595422;
assign addr[8204]= -107043224;
assign addr[8205]= -183355234;
assign addr[8206]= -259434643;
assign addr[8207]= -335184940;
assign addr[8208]= -410510029;
assign addr[8209]= -485314355;
assign addr[8210]= -559503022;
assign addr[8211]= -632981917;
assign addr[8212]= -705657826;
assign addr[8213]= -777438554;
assign addr[8214]= -848233042;
assign addr[8215]= -917951481;
assign addr[8216]= -986505429;
assign addr[8217]= -1053807919;
assign addr[8218]= -1119773573;
assign addr[8219]= -1184318708;
assign addr[8220]= -1247361445;
assign addr[8221]= -1308821808;
assign addr[8222]= -1368621831;
assign addr[8223]= -1426685652;
assign addr[8224]= -1482939614;
assign addr[8225]= -1537312353;
assign addr[8226]= -1589734894;
assign addr[8227]= -1640140734;
assign addr[8228]= -1688465931;
assign addr[8229]= -1734649179;
assign addr[8230]= -1778631892;
assign addr[8231]= -1820358275;
assign addr[8232]= -1859775393;
assign addr[8233]= -1896833245;
assign addr[8234]= -1931484818;
assign addr[8235]= -1963686155;
assign addr[8236]= -1993396407;
assign addr[8237]= -2020577882;
assign addr[8238]= -2045196100;
assign addr[8239]= -2067219829;
assign addr[8240]= -2086621133;
assign addr[8241]= -2103375398;
assign addr[8242]= -2117461370;
assign addr[8243]= -2128861181;
assign addr[8244]= -2137560369;
assign addr[8245]= -2143547897;
assign addr[8246]= -2146816171;
assign addr[8247]= -2147361045;
assign addr[8248]= -2145181827;
assign addr[8249]= -2140281282;
assign addr[8250]= -2132665626;
assign addr[8251]= -2122344521;
assign addr[8252]= -2109331059;
assign addr[8253]= -2093641749;
assign addr[8254]= -2075296495;
assign addr[8255]= -2054318569;
assign addr[8256]= -2030734582;
assign addr[8257]= -2004574453;
assign addr[8258]= -1975871368;
assign addr[8259]= -1944661739;
assign addr[8260]= -1910985158;
assign addr[8261]= -1874884346;
assign addr[8262]= -1836405100;
assign addr[8263]= -1795596234;
assign addr[8264]= -1752509516;
assign addr[8265]= -1707199606;
assign addr[8266]= -1659723983;
assign addr[8267]= -1610142873;
assign addr[8268]= -1558519173;
assign addr[8269]= -1504918373;
assign addr[8270]= -1449408469;
assign addr[8271]= -1392059879;
assign addr[8272]= -1332945355;
assign addr[8273]= -1272139887;
assign addr[8274]= -1209720613;
assign addr[8275]= -1145766716;
assign addr[8276]= -1080359326;
assign addr[8277]= -1013581418;
assign addr[8278]= -945517704;
assign addr[8279]= -876254528;
assign addr[8280]= -805879757;
assign addr[8281]= -734482665;
assign addr[8282]= -662153826;
assign addr[8283]= -588984994;
assign addr[8284]= -515068990;
assign addr[8285]= -440499581;
assign addr[8286]= -365371365;
assign addr[8287]= -289779648;
assign addr[8288]= -213820322;
assign addr[8289]= -137589750;
assign addr[8290]= -61184634;
assign addr[8291]= 15298099;
assign addr[8292]= 91761426;
assign addr[8293]= 168108346;
assign addr[8294]= 244242007;
assign addr[8295]= 320065829;
assign addr[8296]= 395483624;
assign addr[8297]= 470399716;
assign addr[8298]= 544719071;
assign addr[8299]= 618347408;
assign addr[8300]= 691191324;
assign addr[8301]= 763158411;
assign addr[8302]= 834157373;
assign addr[8303]= 904098143;
assign addr[8304]= 972891995;
assign addr[8305]= 1040451659;
assign addr[8306]= 1106691431;
assign addr[8307]= 1171527280;
assign addr[8308]= 1234876957;
assign addr[8309]= 1296660098;
assign addr[8310]= 1356798326;
assign addr[8311]= 1415215352;
assign addr[8312]= 1471837070;
assign addr[8313]= 1526591649;
assign addr[8314]= 1579409630;
assign addr[8315]= 1630224009;
assign addr[8316]= 1678970324;
assign addr[8317]= 1725586737;
assign addr[8318]= 1770014111;
assign addr[8319]= 1812196087;
assign addr[8320]= 1852079154;
assign addr[8321]= 1889612716;
assign addr[8322]= 1924749160;
assign addr[8323]= 1957443913;
assign addr[8324]= 1987655498;
assign addr[8325]= 2015345591;
assign addr[8326]= 2040479063;
assign addr[8327]= 2063024031;
assign addr[8328]= 2082951896;
assign addr[8329]= 2100237377;
assign addr[8330]= 2114858546;
assign addr[8331]= 2126796855;
assign addr[8332]= 2136037160;
assign addr[8333]= 2142567738;
assign addr[8334]= 2146380306;
assign addr[8335]= 2147470025;
assign addr[8336]= 2145835515;
assign addr[8337]= 2141478848;
assign addr[8338]= 2134405552;
assign addr[8339]= 2124624598;
assign addr[8340]= 2112148396;
assign addr[8341]= 2096992772;
assign addr[8342]= 2079176953;
assign addr[8343]= 2058723538;
assign addr[8344]= 2035658475;
assign addr[8345]= 2010011024;
assign addr[8346]= 1981813720;
assign addr[8347]= 1951102334;
assign addr[8348]= 1917915825;
assign addr[8349]= 1882296293;
assign addr[8350]= 1844288924;
assign addr[8351]= 1803941934;
assign addr[8352]= 1761306505;
assign addr[8353]= 1716436725;
assign addr[8354]= 1669389513;
assign addr[8355]= 1620224553;
assign addr[8356]= 1569004214;
assign addr[8357]= 1515793473;
assign addr[8358]= 1460659832;
assign addr[8359]= 1403673233;
assign addr[8360]= 1344905966;
assign addr[8361]= 1284432584;
assign addr[8362]= 1222329801;
assign addr[8363]= 1158676398;
assign addr[8364]= 1093553126;
assign addr[8365]= 1027042599;
assign addr[8366]= 959229189;
assign addr[8367]= 890198924;
assign addr[8368]= 820039373;
assign addr[8369]= 748839539;
assign addr[8370]= 676689746;
assign addr[8371]= 603681519;
assign addr[8372]= 529907477;
assign addr[8373]= 455461206;
assign addr[8374]= 380437148;
assign addr[8375]= 304930476;
assign addr[8376]= 229036977;
assign addr[8377]= 152852926;
assign addr[8378]= 76474970;
assign addr[8379]= 0;
assign addr[8380]= -76474970;
assign addr[8381]= -152852926;
assign addr[8382]= -229036977;
assign addr[8383]= -304930476;
assign addr[8384]= -380437148;
assign addr[8385]= -455461206;
assign addr[8386]= -529907477;
assign addr[8387]= -603681519;
assign addr[8388]= -676689746;
assign addr[8389]= -748839539;
assign addr[8390]= -820039373;
assign addr[8391]= -890198924;
assign addr[8392]= -959229189;
assign addr[8393]= -1027042599;
assign addr[8394]= -1093553126;
assign addr[8395]= -1158676398;
assign addr[8396]= -1222329801;
assign addr[8397]= -1284432584;
assign addr[8398]= -1344905966;
assign addr[8399]= -1403673233;
assign addr[8400]= -1460659832;
assign addr[8401]= -1515793473;
assign addr[8402]= -1569004214;
assign addr[8403]= -1620224553;
assign addr[8404]= -1669389513;
assign addr[8405]= -1716436725;
assign addr[8406]= -1761306505;
assign addr[8407]= -1803941934;
assign addr[8408]= -1844288924;
assign addr[8409]= -1882296293;
assign addr[8410]= -1917915825;
assign addr[8411]= -1951102334;
assign addr[8412]= -1981813720;
assign addr[8413]= -2010011024;
assign addr[8414]= -2035658475;
assign addr[8415]= -2058723538;
assign addr[8416]= -2079176953;
assign addr[8417]= -2096992772;
assign addr[8418]= -2112148396;
assign addr[8419]= -2124624598;
assign addr[8420]= -2134405552;
assign addr[8421]= -2141478848;
assign addr[8422]= -2145835515;
assign addr[8423]= -2147470025;
assign addr[8424]= -2146380306;
assign addr[8425]= -2142567738;
assign addr[8426]= -2136037160;
assign addr[8427]= -2126796855;
assign addr[8428]= -2114858546;
assign addr[8429]= -2100237377;
assign addr[8430]= -2082951896;
assign addr[8431]= -2063024031;
assign addr[8432]= -2040479063;
assign addr[8433]= -2015345591;
assign addr[8434]= -1987655498;
assign addr[8435]= -1957443913;
assign addr[8436]= -1924749160;
assign addr[8437]= -1889612716;
assign addr[8438]= -1852079154;
assign addr[8439]= -1812196087;
assign addr[8440]= -1770014111;
assign addr[8441]= -1725586737;
assign addr[8442]= -1678970324;
assign addr[8443]= -1630224009;
assign addr[8444]= -1579409630;
assign addr[8445]= -1526591649;
assign addr[8446]= -1471837070;
assign addr[8447]= -1415215352;
assign addr[8448]= -1356798326;
assign addr[8449]= -1296660098;
assign addr[8450]= -1234876957;
assign addr[8451]= -1171527280;
assign addr[8452]= -1106691431;
assign addr[8453]= -1040451659;
assign addr[8454]= -972891995;
assign addr[8455]= -904098143;
assign addr[8456]= -834157373;
assign addr[8457]= -763158411;
assign addr[8458]= -691191324;
assign addr[8459]= -618347408;
assign addr[8460]= -544719071;
assign addr[8461]= -470399716;
assign addr[8462]= -395483624;
assign addr[8463]= -320065829;
assign addr[8464]= -244242007;
assign addr[8465]= -168108346;
assign addr[8466]= -91761426;
assign addr[8467]= -15298099;
assign addr[8468]= 61184634;
assign addr[8469]= 137589750;
assign addr[8470]= 213820322;
assign addr[8471]= 289779648;
assign addr[8472]= 365371365;
assign addr[8473]= 440499581;
assign addr[8474]= 515068990;
assign addr[8475]= 588984994;
assign addr[8476]= 662153826;
assign addr[8477]= 734482665;
assign addr[8478]= 805879757;
assign addr[8479]= 876254528;
assign addr[8480]= 945517704;
assign addr[8481]= 1013581418;
assign addr[8482]= 1080359326;
assign addr[8483]= 1145766716;
assign addr[8484]= 1209720613;
assign addr[8485]= 1272139887;
assign addr[8486]= 1332945355;
assign addr[8487]= 1392059879;
assign addr[8488]= 1449408469;
assign addr[8489]= 1504918373;
assign addr[8490]= 1558519173;
assign addr[8491]= 1610142873;
assign addr[8492]= 1659723983;
assign addr[8493]= 1707199606;
assign addr[8494]= 1752509516;
assign addr[8495]= 1795596234;
assign addr[8496]= 1836405100;
assign addr[8497]= 1874884346;
assign addr[8498]= 1910985158;
assign addr[8499]= 1944661739;
assign addr[8500]= 1975871368;
assign addr[8501]= 2004574453;
assign addr[8502]= 2030734582;
assign addr[8503]= 2054318569;
assign addr[8504]= 2075296495;
assign addr[8505]= 2093641749;
assign addr[8506]= 2109331059;
assign addr[8507]= 2122344521;
assign addr[8508]= 2132665626;
assign addr[8509]= 2140281282;
assign addr[8510]= 2145181827;
assign addr[8511]= 2147361045;
assign addr[8512]= 2146816171;
assign addr[8513]= 2143547897;
assign addr[8514]= 2137560369;
assign addr[8515]= 2128861181;
assign addr[8516]= 2117461370;
assign addr[8517]= 2103375398;
assign addr[8518]= 2086621133;
assign addr[8519]= 2067219829;
assign addr[8520]= 2045196100;
assign addr[8521]= 2020577882;
assign addr[8522]= 1993396407;
assign addr[8523]= 1963686155;
assign addr[8524]= 1931484818;
assign addr[8525]= 1896833245;
assign addr[8526]= 1859775393;
assign addr[8527]= 1820358275;
assign addr[8528]= 1778631892;
assign addr[8529]= 1734649179;
assign addr[8530]= 1688465931;
assign addr[8531]= 1640140734;
assign addr[8532]= 1589734894;
assign addr[8533]= 1537312353;
assign addr[8534]= 1482939614;
assign addr[8535]= 1426685652;
assign addr[8536]= 1368621831;
assign addr[8537]= 1308821808;
assign addr[8538]= 1247361445;
assign addr[8539]= 1184318708;
assign addr[8540]= 1119773573;
assign addr[8541]= 1053807919;
assign addr[8542]= 986505429;
assign addr[8543]= 917951481;
assign addr[8544]= 848233042;
assign addr[8545]= 777438554;
assign addr[8546]= 705657826;
assign addr[8547]= 632981917;
assign addr[8548]= 559503022;
assign addr[8549]= 485314355;
assign addr[8550]= 410510029;
assign addr[8551]= 335184940;
assign addr[8552]= 259434643;
assign addr[8553]= 183355234;
assign addr[8554]= 107043224;
assign addr[8555]= 30595422;
assign addr[8556]= -45891193;
assign addr[8557]= -122319591;
assign addr[8558]= -198592817;
assign addr[8559]= -274614114;
assign addr[8560]= -350287041;
assign addr[8561]= -425515602;
assign addr[8562]= -500204365;
assign addr[8563]= -574258580;
assign addr[8564]= -647584304;
assign addr[8565]= -720088517;
assign addr[8566]= -791679244;
assign addr[8567]= -862265664;
assign addr[8568]= -931758235;
assign addr[8569]= -1000068799;
assign addr[8570]= -1067110699;
assign addr[8571]= -1132798888;
assign addr[8572]= -1197050035;
assign addr[8573]= -1259782632;
assign addr[8574]= -1320917099;
assign addr[8575]= -1380375881;
assign addr[8576]= -1438083551;
assign addr[8577]= -1493966902;
assign addr[8578]= -1547955041;
assign addr[8579]= -1599979481;
assign addr[8580]= -1649974225;
assign addr[8581]= -1697875851;
assign addr[8582]= -1743623590;
assign addr[8583]= -1787159411;
assign addr[8584]= -1828428082;
assign addr[8585]= -1867377253;
assign addr[8586]= -1903957513;
assign addr[8587]= -1938122457;
assign addr[8588]= -1969828744;
assign addr[8589]= -1999036154;
assign addr[8590]= -2025707632;
assign addr[8591]= -2049809346;
assign addr[8592]= -2071310720;
assign addr[8593]= -2090184478;
assign addr[8594]= -2106406677;
assign addr[8595]= -2119956737;
assign addr[8596]= -2130817471;
assign addr[8597]= -2138975100;
assign addr[8598]= -2144419275;
assign addr[8599]= -2147143090;
assign addr[8600]= -2147143090;
assign addr[8601]= -2144419275;
assign addr[8602]= -2138975100;
assign addr[8603]= -2130817471;
assign addr[8604]= -2119956737;
assign addr[8605]= -2106406677;
assign addr[8606]= -2090184478;
assign addr[8607]= -2071310720;
assign addr[8608]= -2049809346;
assign addr[8609]= -2025707632;
assign addr[8610]= -1999036154;
assign addr[8611]= -1969828744;
assign addr[8612]= -1938122457;
assign addr[8613]= -1903957513;
assign addr[8614]= -1867377253;
assign addr[8615]= -1828428082;
assign addr[8616]= -1787159411;
assign addr[8617]= -1743623590;
assign addr[8618]= -1697875851;
assign addr[8619]= -1649974225;
assign addr[8620]= -1599979481;
assign addr[8621]= -1547955041;
assign addr[8622]= -1493966902;
assign addr[8623]= -1438083551;
assign addr[8624]= -1380375881;
assign addr[8625]= -1320917099;
assign addr[8626]= -1259782632;
assign addr[8627]= -1197050035;
assign addr[8628]= -1132798888;
assign addr[8629]= -1067110699;
assign addr[8630]= -1000068799;
assign addr[8631]= -931758235;
assign addr[8632]= -862265664;
assign addr[8633]= -791679244;
assign addr[8634]= -720088517;
assign addr[8635]= -647584304;
assign addr[8636]= -574258580;
assign addr[8637]= -500204365;
assign addr[8638]= -425515602;
assign addr[8639]= -350287041;
assign addr[8640]= -274614114;
assign addr[8641]= -198592817;
assign addr[8642]= -122319591;
assign addr[8643]= -45891193;
assign addr[8644]= 30595422;
assign addr[8645]= 107043224;
assign addr[8646]= 183355234;
assign addr[8647]= 259434643;
assign addr[8648]= 335184940;
assign addr[8649]= 410510029;
assign addr[8650]= 485314355;
assign addr[8651]= 559503022;
assign addr[8652]= 632981917;
assign addr[8653]= 705657826;
assign addr[8654]= 777438554;
assign addr[8655]= 848233042;
assign addr[8656]= 917951481;
assign addr[8657]= 986505429;
assign addr[8658]= 1053807919;
assign addr[8659]= 1119773573;
assign addr[8660]= 1184318708;
assign addr[8661]= 1247361445;
assign addr[8662]= 1308821808;
assign addr[8663]= 1368621831;
assign addr[8664]= 1426685652;
assign addr[8665]= 1482939614;
assign addr[8666]= 1537312353;
assign addr[8667]= 1589734894;
assign addr[8668]= 1640140734;
assign addr[8669]= 1688465931;
assign addr[8670]= 1734649179;
assign addr[8671]= 1778631892;
assign addr[8672]= 1820358275;
assign addr[8673]= 1859775393;
assign addr[8674]= 1896833245;
assign addr[8675]= 1931484818;
assign addr[8676]= 1963686155;
assign addr[8677]= 1993396407;
assign addr[8678]= 2020577882;
assign addr[8679]= 2045196100;
assign addr[8680]= 2067219829;
assign addr[8681]= 2086621133;
assign addr[8682]= 2103375398;
assign addr[8683]= 2117461370;
assign addr[8684]= 2128861181;
assign addr[8685]= 2137560369;
assign addr[8686]= 2143547897;
assign addr[8687]= 2146816171;
assign addr[8688]= 2147361045;
assign addr[8689]= 2145181827;
assign addr[8690]= 2140281282;
assign addr[8691]= 2132665626;
assign addr[8692]= 2122344521;
assign addr[8693]= 2109331059;
assign addr[8694]= 2093641749;
assign addr[8695]= 2075296495;
assign addr[8696]= 2054318569;
assign addr[8697]= 2030734582;
assign addr[8698]= 2004574453;
assign addr[8699]= 1975871368;
assign addr[8700]= 1944661739;
assign addr[8701]= 1910985158;
assign addr[8702]= 1874884346;
assign addr[8703]= 1836405100;
assign addr[8704]= 1795596234;
assign addr[8705]= 1752509516;
assign addr[8706]= 1707199606;
assign addr[8707]= 1659723983;
assign addr[8708]= 1610142873;
assign addr[8709]= 1558519173;
assign addr[8710]= 1504918373;
assign addr[8711]= 1449408469;
assign addr[8712]= 1392059879;
assign addr[8713]= 1332945355;
assign addr[8714]= 1272139887;
assign addr[8715]= 1209720613;
assign addr[8716]= 1145766716;
assign addr[8717]= 1080359326;
assign addr[8718]= 1013581418;
assign addr[8719]= 945517704;
assign addr[8720]= 876254528;
assign addr[8721]= 805879757;
assign addr[8722]= 734482665;
assign addr[8723]= 662153826;
assign addr[8724]= 588984994;
assign addr[8725]= 515068990;
assign addr[8726]= 440499581;
assign addr[8727]= 365371365;
assign addr[8728]= 289779648;
assign addr[8729]= 213820322;
assign addr[8730]= 137589750;
assign addr[8731]= 61184634;
assign addr[8732]= -15298099;
assign addr[8733]= -91761426;
assign addr[8734]= -168108346;
assign addr[8735]= -244242007;
assign addr[8736]= -320065829;
assign addr[8737]= -395483624;
assign addr[8738]= -470399716;
assign addr[8739]= -544719071;
assign addr[8740]= -618347408;
assign addr[8741]= -691191324;
assign addr[8742]= -763158411;
assign addr[8743]= -834157373;
assign addr[8744]= -904098143;
assign addr[8745]= -972891995;
assign addr[8746]= -1040451659;
assign addr[8747]= -1106691431;
assign addr[8748]= -1171527280;
assign addr[8749]= -1234876957;
assign addr[8750]= -1296660098;
assign addr[8751]= -1356798326;
assign addr[8752]= -1415215352;
assign addr[8753]= -1471837070;
assign addr[8754]= -1526591649;
assign addr[8755]= -1579409630;
assign addr[8756]= -1630224009;
assign addr[8757]= -1678970324;
assign addr[8758]= -1725586737;
assign addr[8759]= -1770014111;
assign addr[8760]= -1812196087;
assign addr[8761]= -1852079154;
assign addr[8762]= -1889612716;
assign addr[8763]= -1924749160;
assign addr[8764]= -1957443913;
assign addr[8765]= -1987655498;
assign addr[8766]= -2015345591;
assign addr[8767]= -2040479063;
assign addr[8768]= -2063024031;
assign addr[8769]= -2082951896;
assign addr[8770]= -2100237377;
assign addr[8771]= -2114858546;
assign addr[8772]= -2126796855;
assign addr[8773]= -2136037160;
assign addr[8774]= -2142567738;
assign addr[8775]= -2146380306;
assign addr[8776]= -2147470025;
assign addr[8777]= -2145835515;
assign addr[8778]= -2141478848;
assign addr[8779]= -2134405552;
assign addr[8780]= -2124624598;
assign addr[8781]= -2112148396;
assign addr[8782]= -2096992772;
assign addr[8783]= -2079176953;
assign addr[8784]= -2058723538;
assign addr[8785]= -2035658475;
assign addr[8786]= -2010011024;
assign addr[8787]= -1981813720;
assign addr[8788]= -1951102334;
assign addr[8789]= -1917915825;
assign addr[8790]= -1882296293;
assign addr[8791]= -1844288924;
assign addr[8792]= -1803941934;
assign addr[8793]= -1761306505;
assign addr[8794]= -1716436725;
assign addr[8795]= -1669389513;
assign addr[8796]= -1620224553;
assign addr[8797]= -1569004214;
assign addr[8798]= -1515793473;
assign addr[8799]= -1460659832;
assign addr[8800]= -1403673233;
assign addr[8801]= -1344905966;
assign addr[8802]= -1284432584;
assign addr[8803]= -1222329801;
assign addr[8804]= -1158676398;
assign addr[8805]= -1093553126;
assign addr[8806]= -1027042599;
assign addr[8807]= -959229189;
assign addr[8808]= -890198924;
assign addr[8809]= -820039373;
assign addr[8810]= -748839539;
assign addr[8811]= -676689746;
assign addr[8812]= -603681519;
assign addr[8813]= -529907477;
assign addr[8814]= -455461206;
assign addr[8815]= -380437148;
assign addr[8816]= -304930476;
assign addr[8817]= -229036977;
assign addr[8818]= -152852926;
assign addr[8819]= -76474970;
assign addr[8820]= 0;
assign addr[8821]= 76474970;
assign addr[8822]= 152852926;
assign addr[8823]= 229036977;
assign addr[8824]= 304930476;
assign addr[8825]= 380437148;
assign addr[8826]= 455461206;
assign addr[8827]= 529907477;
assign addr[8828]= 603681519;
assign addr[8829]= 676689746;
assign addr[8830]= 748839539;
assign addr[8831]= 820039373;
assign addr[8832]= 890198924;
assign addr[8833]= 959229189;
assign addr[8834]= 1027042599;
assign addr[8835]= 1093553126;
assign addr[8836]= 1158676398;
assign addr[8837]= 1222329801;
assign addr[8838]= 1284432584;
assign addr[8839]= 1344905966;
assign addr[8840]= 1403673233;
assign addr[8841]= 1460659832;
assign addr[8842]= 1515793473;
assign addr[8843]= 1569004214;
assign addr[8844]= 1620224553;
assign addr[8845]= 1669389513;
assign addr[8846]= 1716436725;
assign addr[8847]= 1761306505;
assign addr[8848]= 1803941934;
assign addr[8849]= 1844288924;
assign addr[8850]= 1882296293;
assign addr[8851]= 1917915825;
assign addr[8852]= 1951102334;
assign addr[8853]= 1981813720;
assign addr[8854]= 2010011024;
assign addr[8855]= 2035658475;
assign addr[8856]= 2058723538;
assign addr[8857]= 2079176953;
assign addr[8858]= 2096992772;
assign addr[8859]= 2112148396;
assign addr[8860]= 2124624598;
assign addr[8861]= 2134405552;
assign addr[8862]= 2141478848;
assign addr[8863]= 2145835515;
assign addr[8864]= 2147470025;
assign addr[8865]= 2146380306;
assign addr[8866]= 2142567738;
assign addr[8867]= 2136037160;
assign addr[8868]= 2126796855;
assign addr[8869]= 2114858546;
assign addr[8870]= 2100237377;
assign addr[8871]= 2082951896;
assign addr[8872]= 2063024031;
assign addr[8873]= 2040479063;
assign addr[8874]= 2015345591;
assign addr[8875]= 1987655498;
assign addr[8876]= 1957443913;
assign addr[8877]= 1924749160;
assign addr[8878]= 1889612716;
assign addr[8879]= 1852079154;
assign addr[8880]= 1812196087;
assign addr[8881]= 1770014111;
assign addr[8882]= 1725586737;
assign addr[8883]= 1678970324;
assign addr[8884]= 1630224009;
assign addr[8885]= 1579409630;
assign addr[8886]= 1526591649;
assign addr[8887]= 1471837070;
assign addr[8888]= 1415215352;
assign addr[8889]= 1356798326;
assign addr[8890]= 1296660098;
assign addr[8891]= 1234876957;
assign addr[8892]= 1171527280;
assign addr[8893]= 1106691431;
assign addr[8894]= 1040451659;
assign addr[8895]= 972891995;
assign addr[8896]= 904098143;
assign addr[8897]= 834157373;
assign addr[8898]= 763158411;
assign addr[8899]= 691191324;
assign addr[8900]= 618347408;
assign addr[8901]= 544719071;
assign addr[8902]= 470399716;
assign addr[8903]= 395483624;
assign addr[8904]= 320065829;
assign addr[8905]= 244242007;
assign addr[8906]= 168108346;
assign addr[8907]= 91761426;
assign addr[8908]= 15298099;
assign addr[8909]= -61184634;
assign addr[8910]= -137589750;
assign addr[8911]= -213820322;
assign addr[8912]= -289779648;
assign addr[8913]= -365371365;
assign addr[8914]= -440499581;
assign addr[8915]= -515068990;
assign addr[8916]= -588984994;
assign addr[8917]= -662153826;
assign addr[8918]= -734482665;
assign addr[8919]= -805879757;
assign addr[8920]= -876254528;
assign addr[8921]= -945517704;
assign addr[8922]= -1013581418;
assign addr[8923]= -1080359326;
assign addr[8924]= -1145766716;
assign addr[8925]= -1209720613;
assign addr[8926]= -1272139887;
assign addr[8927]= -1332945355;
assign addr[8928]= -1392059879;
assign addr[8929]= -1449408469;
assign addr[8930]= -1504918373;
assign addr[8931]= -1558519173;
assign addr[8932]= -1610142873;
assign addr[8933]= -1659723983;
assign addr[8934]= -1707199606;
assign addr[8935]= -1752509516;
assign addr[8936]= -1795596234;
assign addr[8937]= -1836405100;
assign addr[8938]= -1874884346;
assign addr[8939]= -1910985158;
assign addr[8940]= -1944661739;
assign addr[8941]= -1975871368;
assign addr[8942]= -2004574453;
assign addr[8943]= -2030734582;
assign addr[8944]= -2054318569;
assign addr[8945]= -2075296495;
assign addr[8946]= -2093641749;
assign addr[8947]= -2109331059;
assign addr[8948]= -2122344521;
assign addr[8949]= -2132665626;
assign addr[8950]= -2140281282;
assign addr[8951]= -2145181827;
assign addr[8952]= -2147361045;
assign addr[8953]= -2146816171;
assign addr[8954]= -2143547897;
assign addr[8955]= -2137560369;
assign addr[8956]= -2128861181;
assign addr[8957]= -2117461370;
assign addr[8958]= -2103375398;
assign addr[8959]= -2086621133;
assign addr[8960]= -2067219829;
assign addr[8961]= -2045196100;
assign addr[8962]= -2020577882;
assign addr[8963]= -1993396407;
assign addr[8964]= -1963686155;
assign addr[8965]= -1931484818;
assign addr[8966]= -1896833245;
assign addr[8967]= -1859775393;
assign addr[8968]= -1820358275;
assign addr[8969]= -1778631892;
assign addr[8970]= -1734649179;
assign addr[8971]= -1688465931;
assign addr[8972]= -1640140734;
assign addr[8973]= -1589734894;
assign addr[8974]= -1537312353;
assign addr[8975]= -1482939614;
assign addr[8976]= -1426685652;
assign addr[8977]= -1368621831;
assign addr[8978]= -1308821808;
assign addr[8979]= -1247361445;
assign addr[8980]= -1184318708;
assign addr[8981]= -1119773573;
assign addr[8982]= -1053807919;
assign addr[8983]= -986505429;
assign addr[8984]= -917951481;
assign addr[8985]= -848233042;
assign addr[8986]= -777438554;
assign addr[8987]= -705657826;
assign addr[8988]= -632981917;
assign addr[8989]= -559503022;
assign addr[8990]= -485314355;
assign addr[8991]= -410510029;
assign addr[8992]= -335184940;
assign addr[8993]= -259434643;
assign addr[8994]= -183355234;
assign addr[8995]= -107043224;
assign addr[8996]= -30595422;
assign addr[8997]= 45891193;
assign addr[8998]= 122319591;
assign addr[8999]= 198592817;
assign addr[9000]= 274614114;
assign addr[9001]= 350287041;
assign addr[9002]= 425515602;
assign addr[9003]= 500204365;
assign addr[9004]= 574258580;
assign addr[9005]= 647584304;
assign addr[9006]= 720088517;
assign addr[9007]= 791679244;
assign addr[9008]= 862265664;
assign addr[9009]= 931758235;
assign addr[9010]= 1000068799;
assign addr[9011]= 1067110699;
assign addr[9012]= 1132798888;
assign addr[9013]= 1197050035;
assign addr[9014]= 1259782632;
assign addr[9015]= 1320917099;
assign addr[9016]= 1380375881;
assign addr[9017]= 1438083551;
assign addr[9018]= 1493966902;
assign addr[9019]= 1547955041;
assign addr[9020]= 1599979481;
assign addr[9021]= 1649974225;
assign addr[9022]= 1697875851;
assign addr[9023]= 1743623590;
assign addr[9024]= 1787159411;
assign addr[9025]= 1828428082;
assign addr[9026]= 1867377253;
assign addr[9027]= 1903957513;
assign addr[9028]= 1938122457;
assign addr[9029]= 1969828744;
assign addr[9030]= 1999036154;
assign addr[9031]= 2025707632;
assign addr[9032]= 2049809346;
assign addr[9033]= 2071310720;
assign addr[9034]= 2090184478;
assign addr[9035]= 2106406677;
assign addr[9036]= 2119956737;
assign addr[9037]= 2130817471;
assign addr[9038]= 2138975100;
assign addr[9039]= 2144419275;
assign addr[9040]= 2147143090;
assign addr[9041]= 2147143090;
assign addr[9042]= 2144419275;
assign addr[9043]= 2138975100;
assign addr[9044]= 2130817471;
assign addr[9045]= 2119956737;
assign addr[9046]= 2106406677;
assign addr[9047]= 2090184478;
assign addr[9048]= 2071310720;
assign addr[9049]= 2049809346;
assign addr[9050]= 2025707632;
assign addr[9051]= 1999036154;
assign addr[9052]= 1969828744;
assign addr[9053]= 1938122457;
assign addr[9054]= 1903957513;
assign addr[9055]= 1867377253;
assign addr[9056]= 1828428082;
assign addr[9057]= 1787159411;
assign addr[9058]= 1743623590;
assign addr[9059]= 1697875851;
assign addr[9060]= 1649974225;
assign addr[9061]= 1599979481;
assign addr[9062]= 1547955041;
assign addr[9063]= 1493966902;
assign addr[9064]= 1438083551;
assign addr[9065]= 1380375881;
assign addr[9066]= 1320917099;
assign addr[9067]= 1259782632;
assign addr[9068]= 1197050035;
assign addr[9069]= 1132798888;
assign addr[9070]= 1067110699;
assign addr[9071]= 1000068799;
assign addr[9072]= 931758235;
assign addr[9073]= 862265664;
assign addr[9074]= 791679244;
assign addr[9075]= 720088517;
assign addr[9076]= 647584304;
assign addr[9077]= 574258580;
assign addr[9078]= 500204365;
assign addr[9079]= 425515602;
assign addr[9080]= 350287041;
assign addr[9081]= 274614114;
assign addr[9082]= 198592817;
assign addr[9083]= 122319591;
assign addr[9084]= 45891193;
assign addr[9085]= -30595422;
assign addr[9086]= -107043224;
assign addr[9087]= -183355234;
assign addr[9088]= -259434643;
assign addr[9089]= -335184940;
assign addr[9090]= -410510029;
assign addr[9091]= -485314355;
assign addr[9092]= -559503022;
assign addr[9093]= -632981917;
assign addr[9094]= -705657826;
assign addr[9095]= -777438554;
assign addr[9096]= -848233042;
assign addr[9097]= -917951481;
assign addr[9098]= -986505429;
assign addr[9099]= -1053807919;
assign addr[9100]= -1119773573;
assign addr[9101]= -1184318708;
assign addr[9102]= -1247361445;
assign addr[9103]= -1308821808;
assign addr[9104]= -1368621831;
assign addr[9105]= -1426685652;
assign addr[9106]= -1482939614;
assign addr[9107]= -1537312353;
assign addr[9108]= -1589734894;
assign addr[9109]= -1640140734;
assign addr[9110]= -1688465931;
assign addr[9111]= -1734649179;
assign addr[9112]= -1778631892;
assign addr[9113]= -1820358275;
assign addr[9114]= -1859775393;
assign addr[9115]= -1896833245;
assign addr[9116]= -1931484818;
assign addr[9117]= -1963686155;
assign addr[9118]= -1993396407;
assign addr[9119]= -2020577882;
assign addr[9120]= -2045196100;
assign addr[9121]= -2067219829;
assign addr[9122]= -2086621133;
assign addr[9123]= -2103375398;
assign addr[9124]= -2117461370;
assign addr[9125]= -2128861181;
assign addr[9126]= -2137560369;
assign addr[9127]= -2143547897;
assign addr[9128]= -2146816171;
assign addr[9129]= -2147361045;
assign addr[9130]= -2145181827;
assign addr[9131]= -2140281282;
assign addr[9132]= -2132665626;
assign addr[9133]= -2122344521;
assign addr[9134]= -2109331059;
assign addr[9135]= -2093641749;
assign addr[9136]= -2075296495;
assign addr[9137]= -2054318569;
assign addr[9138]= -2030734582;
assign addr[9139]= -2004574453;
assign addr[9140]= -1975871368;
assign addr[9141]= -1944661739;
assign addr[9142]= -1910985158;
assign addr[9143]= -1874884346;
assign addr[9144]= -1836405100;
assign addr[9145]= -1795596234;
assign addr[9146]= -1752509516;
assign addr[9147]= -1707199606;
assign addr[9148]= -1659723983;
assign addr[9149]= -1610142873;
assign addr[9150]= -1558519173;
assign addr[9151]= -1504918373;
assign addr[9152]= -1449408469;
assign addr[9153]= -1392059879;
assign addr[9154]= -1332945355;
assign addr[9155]= -1272139887;
assign addr[9156]= -1209720613;
assign addr[9157]= -1145766716;
assign addr[9158]= -1080359326;
assign addr[9159]= -1013581418;
assign addr[9160]= -945517704;
assign addr[9161]= -876254528;
assign addr[9162]= -805879757;
assign addr[9163]= -734482665;
assign addr[9164]= -662153826;
assign addr[9165]= -588984994;
assign addr[9166]= -515068990;
assign addr[9167]= -440499581;
assign addr[9168]= -365371365;
assign addr[9169]= -289779648;
assign addr[9170]= -213820322;
assign addr[9171]= -137589750;
assign addr[9172]= -61184634;
assign addr[9173]= 15298099;
assign addr[9174]= 91761426;
assign addr[9175]= 168108346;
assign addr[9176]= 244242007;
assign addr[9177]= 320065829;
assign addr[9178]= 395483624;
assign addr[9179]= 470399716;
assign addr[9180]= 544719071;
assign addr[9181]= 618347408;
assign addr[9182]= 691191324;
assign addr[9183]= 763158411;
assign addr[9184]= 834157373;
assign addr[9185]= 904098143;
assign addr[9186]= 972891995;
assign addr[9187]= 1040451659;
assign addr[9188]= 1106691431;
assign addr[9189]= 1171527280;
assign addr[9190]= 1234876957;
assign addr[9191]= 1296660098;
assign addr[9192]= 1356798326;
assign addr[9193]= 1415215352;
assign addr[9194]= 1471837070;
assign addr[9195]= 1526591649;
assign addr[9196]= 1579409630;
assign addr[9197]= 1630224009;
assign addr[9198]= 1678970324;
assign addr[9199]= 1725586737;
assign addr[9200]= 1770014111;
assign addr[9201]= 1812196087;
assign addr[9202]= 1852079154;
assign addr[9203]= 1889612716;
assign addr[9204]= 1924749160;
assign addr[9205]= 1957443913;
assign addr[9206]= 1987655498;
assign addr[9207]= 2015345591;
assign addr[9208]= 2040479063;
assign addr[9209]= 2063024031;
assign addr[9210]= 2082951896;
assign addr[9211]= 2100237377;
assign addr[9212]= 2114858546;
assign addr[9213]= 2126796855;
assign addr[9214]= 2136037160;
assign addr[9215]= 2142567738;
assign addr[9216]= 2146380306;
assign addr[9217]= 2147470025;
assign addr[9218]= 2145835515;
assign addr[9219]= 2141478848;
assign addr[9220]= 2134405552;
assign addr[9221]= 2124624598;
assign addr[9222]= 2112148396;
assign addr[9223]= 2096992772;
assign addr[9224]= 2079176953;
assign addr[9225]= 2058723538;
assign addr[9226]= 2035658475;
assign addr[9227]= 2010011024;
assign addr[9228]= 1981813720;
assign addr[9229]= 1951102334;
assign addr[9230]= 1917915825;
assign addr[9231]= 1882296293;
assign addr[9232]= 1844288924;
assign addr[9233]= 1803941934;
assign addr[9234]= 1761306505;
assign addr[9235]= 1716436725;
assign addr[9236]= 1669389513;
assign addr[9237]= 1620224553;
assign addr[9238]= 1569004214;
assign addr[9239]= 1515793473;
assign addr[9240]= 1460659832;
assign addr[9241]= 1403673233;
assign addr[9242]= 1344905966;
assign addr[9243]= 1284432584;
assign addr[9244]= 1222329801;
assign addr[9245]= 1158676398;
assign addr[9246]= 1093553126;
assign addr[9247]= 1027042599;
assign addr[9248]= 959229189;
assign addr[9249]= 890198924;
assign addr[9250]= 820039373;
assign addr[9251]= 748839539;
assign addr[9252]= 676689746;
assign addr[9253]= 603681519;
assign addr[9254]= 529907477;
assign addr[9255]= 455461206;
assign addr[9256]= 380437148;
assign addr[9257]= 304930476;
assign addr[9258]= 229036977;
assign addr[9259]= 152852926;
assign addr[9260]= 76474970;
assign addr[9261]= 0;
assign addr[9262]= -76474970;
assign addr[9263]= -152852926;
assign addr[9264]= -229036977;
assign addr[9265]= -304930476;
assign addr[9266]= -380437148;
assign addr[9267]= -455461206;
assign addr[9268]= -529907477;
assign addr[9269]= -603681519;
assign addr[9270]= -676689746;
assign addr[9271]= -748839539;
assign addr[9272]= -820039373;
assign addr[9273]= -890198924;
assign addr[9274]= -959229189;
assign addr[9275]= -1027042599;
assign addr[9276]= -1093553126;
assign addr[9277]= -1158676398;
assign addr[9278]= -1222329801;
assign addr[9279]= -1284432584;
assign addr[9280]= -1344905966;
assign addr[9281]= -1403673233;
assign addr[9282]= -1460659832;
assign addr[9283]= -1515793473;
assign addr[9284]= -1569004214;
assign addr[9285]= -1620224553;
assign addr[9286]= -1669389513;
assign addr[9287]= -1716436725;
assign addr[9288]= -1761306505;
assign addr[9289]= -1803941934;
assign addr[9290]= -1844288924;
assign addr[9291]= -1882296293;
assign addr[9292]= -1917915825;
assign addr[9293]= -1951102334;
assign addr[9294]= -1981813720;
assign addr[9295]= -2010011024;
assign addr[9296]= -2035658475;
assign addr[9297]= -2058723538;
assign addr[9298]= -2079176953;
assign addr[9299]= -2096992772;
assign addr[9300]= -2112148396;
assign addr[9301]= -2124624598;
assign addr[9302]= -2134405552;
assign addr[9303]= -2141478848;
assign addr[9304]= -2145835515;
assign addr[9305]= -2147470025;
assign addr[9306]= -2146380306;
assign addr[9307]= -2142567738;
assign addr[9308]= -2136037160;
assign addr[9309]= -2126796855;
assign addr[9310]= -2114858546;
assign addr[9311]= -2100237377;
assign addr[9312]= -2082951896;
assign addr[9313]= -2063024031;
assign addr[9314]= -2040479063;
assign addr[9315]= -2015345591;
assign addr[9316]= -1987655498;
assign addr[9317]= -1957443913;
assign addr[9318]= -1924749160;
assign addr[9319]= -1889612716;
assign addr[9320]= -1852079154;
assign addr[9321]= -1812196087;
assign addr[9322]= -1770014111;
assign addr[9323]= -1725586737;
assign addr[9324]= -1678970324;
assign addr[9325]= -1630224009;
assign addr[9326]= -1579409630;
assign addr[9327]= -1526591649;
assign addr[9328]= -1471837070;
assign addr[9329]= -1415215352;
assign addr[9330]= -1356798326;
assign addr[9331]= -1296660098;
assign addr[9332]= -1234876957;
assign addr[9333]= -1171527280;
assign addr[9334]= -1106691431;
assign addr[9335]= -1040451659;
assign addr[9336]= -972891995;
assign addr[9337]= -904098143;
assign addr[9338]= -834157373;
assign addr[9339]= -763158411;
assign addr[9340]= -691191324;
assign addr[9341]= -618347408;
assign addr[9342]= -544719071;
assign addr[9343]= -470399716;
assign addr[9344]= -395483624;
assign addr[9345]= -320065829;
assign addr[9346]= -244242007;
assign addr[9347]= -168108346;
assign addr[9348]= -91761426;
assign addr[9349]= -15298099;
assign addr[9350]= 61184634;
assign addr[9351]= 137589750;
assign addr[9352]= 213820322;
assign addr[9353]= 289779648;
assign addr[9354]= 365371365;
assign addr[9355]= 440499581;
assign addr[9356]= 515068990;
assign addr[9357]= 588984994;
assign addr[9358]= 662153826;
assign addr[9359]= 734482665;
assign addr[9360]= 805879757;
assign addr[9361]= 876254528;
assign addr[9362]= 945517704;
assign addr[9363]= 1013581418;
assign addr[9364]= 1080359326;
assign addr[9365]= 1145766716;
assign addr[9366]= 1209720613;
assign addr[9367]= 1272139887;
assign addr[9368]= 1332945355;
assign addr[9369]= 1392059879;
assign addr[9370]= 1449408469;
assign addr[9371]= 1504918373;
assign addr[9372]= 1558519173;
assign addr[9373]= 1610142873;
assign addr[9374]= 1659723983;
assign addr[9375]= 1707199606;
assign addr[9376]= 1752509516;
assign addr[9377]= 1795596234;
assign addr[9378]= 1836405100;
assign addr[9379]= 1874884346;
assign addr[9380]= 1910985158;
assign addr[9381]= 1944661739;
assign addr[9382]= 1975871368;
assign addr[9383]= 2004574453;
assign addr[9384]= 2030734582;
assign addr[9385]= 2054318569;
assign addr[9386]= 2075296495;
assign addr[9387]= 2093641749;
assign addr[9388]= 2109331059;
assign addr[9389]= 2122344521;
assign addr[9390]= 2132665626;
assign addr[9391]= 2140281282;
assign addr[9392]= 2145181827;
assign addr[9393]= 2147361045;
assign addr[9394]= 2146816171;
assign addr[9395]= 2143547897;
assign addr[9396]= 2137560369;
assign addr[9397]= 2128861181;
assign addr[9398]= 2117461370;
assign addr[9399]= 2103375398;
assign addr[9400]= 2086621133;
assign addr[9401]= 2067219829;
assign addr[9402]= 2045196100;
assign addr[9403]= 2020577882;
assign addr[9404]= 1993396407;
assign addr[9405]= 1963686155;
assign addr[9406]= 1931484818;
assign addr[9407]= 1896833245;
assign addr[9408]= 1859775393;
assign addr[9409]= 1820358275;
assign addr[9410]= 1778631892;
assign addr[9411]= 1734649179;
assign addr[9412]= 1688465931;
assign addr[9413]= 1640140734;
assign addr[9414]= 1589734894;
assign addr[9415]= 1537312353;
assign addr[9416]= 1482939614;
assign addr[9417]= 1426685652;
assign addr[9418]= 1368621831;
assign addr[9419]= 1308821808;
assign addr[9420]= 1247361445;
assign addr[9421]= 1184318708;
assign addr[9422]= 1119773573;
assign addr[9423]= 1053807919;
assign addr[9424]= 986505429;
assign addr[9425]= 917951481;
assign addr[9426]= 848233042;
assign addr[9427]= 777438554;
assign addr[9428]= 705657826;
assign addr[9429]= 632981917;
assign addr[9430]= 559503022;
assign addr[9431]= 485314355;
assign addr[9432]= 410510029;
assign addr[9433]= 335184940;
assign addr[9434]= 259434643;
assign addr[9435]= 183355234;
assign addr[9436]= 107043224;
assign addr[9437]= 30595422;
assign addr[9438]= -45891193;
assign addr[9439]= -122319591;
assign addr[9440]= -198592817;
assign addr[9441]= -274614114;
assign addr[9442]= -350287041;
assign addr[9443]= -425515602;
assign addr[9444]= -500204365;
assign addr[9445]= -574258580;
assign addr[9446]= -647584304;
assign addr[9447]= -720088517;
assign addr[9448]= -791679244;
assign addr[9449]= -862265664;
assign addr[9450]= -931758235;
assign addr[9451]= -1000068799;
assign addr[9452]= -1067110699;
assign addr[9453]= -1132798888;
assign addr[9454]= -1197050035;
assign addr[9455]= -1259782632;
assign addr[9456]= -1320917099;
assign addr[9457]= -1380375881;
assign addr[9458]= -1438083551;
assign addr[9459]= -1493966902;
assign addr[9460]= -1547955041;
assign addr[9461]= -1599979481;
assign addr[9462]= -1649974225;
assign addr[9463]= -1697875851;
assign addr[9464]= -1743623590;
assign addr[9465]= -1787159411;
assign addr[9466]= -1828428082;
assign addr[9467]= -1867377253;
assign addr[9468]= -1903957513;
assign addr[9469]= -1938122457;
assign addr[9470]= -1969828744;
assign addr[9471]= -1999036154;
assign addr[9472]= -2025707632;
assign addr[9473]= -2049809346;
assign addr[9474]= -2071310720;
assign addr[9475]= -2090184478;
assign addr[9476]= -2106406677;
assign addr[9477]= -2119956737;
assign addr[9478]= -2130817471;
assign addr[9479]= -2138975100;
assign addr[9480]= -2144419275;
assign addr[9481]= -2147143090;
assign addr[9482]= -2147143090;
assign addr[9483]= -2144419275;
assign addr[9484]= -2138975100;
assign addr[9485]= -2130817471;
assign addr[9486]= -2119956737;
assign addr[9487]= -2106406677;
assign addr[9488]= -2090184478;
assign addr[9489]= -2071310720;
assign addr[9490]= -2049809346;
assign addr[9491]= -2025707632;
assign addr[9492]= -1999036154;
assign addr[9493]= -1969828744;
assign addr[9494]= -1938122457;
assign addr[9495]= -1903957513;
assign addr[9496]= -1867377253;
assign addr[9497]= -1828428082;
assign addr[9498]= -1787159411;
assign addr[9499]= -1743623590;
assign addr[9500]= -1697875851;
assign addr[9501]= -1649974225;
assign addr[9502]= -1599979481;
assign addr[9503]= -1547955041;
assign addr[9504]= -1493966902;
assign addr[9505]= -1438083551;
assign addr[9506]= -1380375881;
assign addr[9507]= -1320917099;
assign addr[9508]= -1259782632;
assign addr[9509]= -1197050035;
assign addr[9510]= -1132798888;
assign addr[9511]= -1067110699;
assign addr[9512]= -1000068799;
assign addr[9513]= -931758235;
assign addr[9514]= -862265664;
assign addr[9515]= -791679244;
assign addr[9516]= -720088517;
assign addr[9517]= -647584304;
assign addr[9518]= -574258580;
assign addr[9519]= -500204365;
assign addr[9520]= -425515602;
assign addr[9521]= -350287041;
assign addr[9522]= -274614114;
assign addr[9523]= -198592817;
assign addr[9524]= -122319591;
assign addr[9525]= -45891193;
assign addr[9526]= 30595422;
assign addr[9527]= 107043224;
assign addr[9528]= 183355234;
assign addr[9529]= 259434643;
assign addr[9530]= 335184940;
assign addr[9531]= 410510029;
assign addr[9532]= 485314355;
assign addr[9533]= 559503022;
assign addr[9534]= 632981917;
assign addr[9535]= 705657826;
assign addr[9536]= 777438554;
assign addr[9537]= 848233042;
assign addr[9538]= 917951481;
assign addr[9539]= 986505429;
assign addr[9540]= 1053807919;
assign addr[9541]= 1119773573;
assign addr[9542]= 1184318708;
assign addr[9543]= 1247361445;
assign addr[9544]= 1308821808;
assign addr[9545]= 1368621831;
assign addr[9546]= 1426685652;
assign addr[9547]= 1482939614;
assign addr[9548]= 1537312353;
assign addr[9549]= 1589734894;
assign addr[9550]= 1640140734;
assign addr[9551]= 1688465931;
assign addr[9552]= 1734649179;
assign addr[9553]= 1778631892;
assign addr[9554]= 1820358275;
assign addr[9555]= 1859775393;
assign addr[9556]= 1896833245;
assign addr[9557]= 1931484818;
assign addr[9558]= 1963686155;
assign addr[9559]= 1993396407;
assign addr[9560]= 2020577882;
assign addr[9561]= 2045196100;
assign addr[9562]= 2067219829;
assign addr[9563]= 2086621133;
assign addr[9564]= 2103375398;
assign addr[9565]= 2117461370;
assign addr[9566]= 2128861181;
assign addr[9567]= 2137560369;
assign addr[9568]= 2143547897;
assign addr[9569]= 2146816171;
assign addr[9570]= 2147361045;
assign addr[9571]= 2145181827;
assign addr[9572]= 2140281282;
assign addr[9573]= 2132665626;
assign addr[9574]= 2122344521;
assign addr[9575]= 2109331059;
assign addr[9576]= 2093641749;
assign addr[9577]= 2075296495;
assign addr[9578]= 2054318569;
assign addr[9579]= 2030734582;
assign addr[9580]= 2004574453;
assign addr[9581]= 1975871368;
assign addr[9582]= 1944661739;
assign addr[9583]= 1910985158;
assign addr[9584]= 1874884346;
assign addr[9585]= 1836405100;
assign addr[9586]= 1795596234;
assign addr[9587]= 1752509516;
assign addr[9588]= 1707199606;
assign addr[9589]= 1659723983;
assign addr[9590]= 1610142873;
assign addr[9591]= 1558519173;
assign addr[9592]= 1504918373;
assign addr[9593]= 1449408469;
assign addr[9594]= 1392059879;
assign addr[9595]= 1332945355;
assign addr[9596]= 1272139887;
assign addr[9597]= 1209720613;
assign addr[9598]= 1145766716;
assign addr[9599]= 1080359326;
assign addr[9600]= 1013581418;
assign addr[9601]= 945517704;
assign addr[9602]= 876254528;
assign addr[9603]= 805879757;
assign addr[9604]= 734482665;
assign addr[9605]= 662153826;
assign addr[9606]= 588984994;
assign addr[9607]= 515068990;
assign addr[9608]= 440499581;
assign addr[9609]= 365371365;
assign addr[9610]= 289779648;
assign addr[9611]= 213820322;
assign addr[9612]= 137589750;
assign addr[9613]= 61184634;
assign addr[9614]= -15298099;
assign addr[9615]= -91761426;
assign addr[9616]= -168108346;
assign addr[9617]= -244242007;
assign addr[9618]= -320065829;
assign addr[9619]= -395483624;
assign addr[9620]= -470399716;
assign addr[9621]= -544719071;
assign addr[9622]= -618347408;
assign addr[9623]= -691191324;
assign addr[9624]= -763158411;
assign addr[9625]= -834157373;
assign addr[9626]= -904098143;
assign addr[9627]= -972891995;
assign addr[9628]= -1040451659;
assign addr[9629]= -1106691431;
assign addr[9630]= -1171527280;
assign addr[9631]= -1234876957;
assign addr[9632]= -1296660098;
assign addr[9633]= -1356798326;
assign addr[9634]= -1415215352;
assign addr[9635]= -1471837070;
assign addr[9636]= -1526591649;
assign addr[9637]= -1579409630;
assign addr[9638]= -1630224009;
assign addr[9639]= -1678970324;
assign addr[9640]= -1725586737;
assign addr[9641]= -1770014111;
assign addr[9642]= -1812196087;
assign addr[9643]= -1852079154;
assign addr[9644]= -1889612716;
assign addr[9645]= -1924749160;
assign addr[9646]= -1957443913;
assign addr[9647]= -1987655498;
assign addr[9648]= -2015345591;
assign addr[9649]= -2040479063;
assign addr[9650]= -2063024031;
assign addr[9651]= -2082951896;
assign addr[9652]= -2100237377;
assign addr[9653]= -2114858546;
assign addr[9654]= -2126796855;
assign addr[9655]= -2136037160;
assign addr[9656]= -2142567738;
assign addr[9657]= -2146380306;
assign addr[9658]= -2147470025;
assign addr[9659]= -2145835515;
assign addr[9660]= -2141478848;
assign addr[9661]= -2134405552;
assign addr[9662]= -2124624598;
assign addr[9663]= -2112148396;
assign addr[9664]= -2096992772;
assign addr[9665]= -2079176953;
assign addr[9666]= -2058723538;
assign addr[9667]= -2035658475;
assign addr[9668]= -2010011024;
assign addr[9669]= -1981813720;
assign addr[9670]= -1951102334;
assign addr[9671]= -1917915825;
assign addr[9672]= -1882296293;
assign addr[9673]= -1844288924;
assign addr[9674]= -1803941934;
assign addr[9675]= -1761306505;
assign addr[9676]= -1716436725;
assign addr[9677]= -1669389513;
assign addr[9678]= -1620224553;
assign addr[9679]= -1569004214;
assign addr[9680]= -1515793473;
assign addr[9681]= -1460659832;
assign addr[9682]= -1403673233;
assign addr[9683]= -1344905966;
assign addr[9684]= -1284432584;
assign addr[9685]= -1222329801;
assign addr[9686]= -1158676398;
assign addr[9687]= -1093553126;
assign addr[9688]= -1027042599;
assign addr[9689]= -959229189;
assign addr[9690]= -890198924;
assign addr[9691]= -820039373;
assign addr[9692]= -748839539;
assign addr[9693]= -676689746;
assign addr[9694]= -603681519;
assign addr[9695]= -529907477;
assign addr[9696]= -455461206;
assign addr[9697]= -380437148;
assign addr[9698]= -304930476;
assign addr[9699]= -229036977;
assign addr[9700]= -152852926;
assign addr[9701]= -76474970;
assign addr[9702]= 0;
assign addr[9703]= 76474970;
assign addr[9704]= 152852926;
assign addr[9705]= 229036977;
assign addr[9706]= 304930476;
assign addr[9707]= 380437148;
assign addr[9708]= 455461206;
assign addr[9709]= 529907477;
assign addr[9710]= 603681519;
assign addr[9711]= 676689746;
assign addr[9712]= 748839539;
assign addr[9713]= 820039373;
assign addr[9714]= 890198924;
assign addr[9715]= 959229189;
assign addr[9716]= 1027042599;
assign addr[9717]= 1093553126;
assign addr[9718]= 1158676398;
assign addr[9719]= 1222329801;
assign addr[9720]= 1284432584;
assign addr[9721]= 1344905966;
assign addr[9722]= 1403673233;
assign addr[9723]= 1460659832;
assign addr[9724]= 1515793473;
assign addr[9725]= 1569004214;
assign addr[9726]= 1620224553;
assign addr[9727]= 1669389513;
assign addr[9728]= 1716436725;
assign addr[9729]= 1761306505;
assign addr[9730]= 1803941934;
assign addr[9731]= 1844288924;
assign addr[9732]= 1882296293;
assign addr[9733]= 1917915825;
assign addr[9734]= 1951102334;
assign addr[9735]= 1981813720;
assign addr[9736]= 2010011024;
assign addr[9737]= 2035658475;
assign addr[9738]= 2058723538;
assign addr[9739]= 2079176953;
assign addr[9740]= 2096992772;
assign addr[9741]= 2112148396;
assign addr[9742]= 2124624598;
assign addr[9743]= 2134405552;
assign addr[9744]= 2141478848;
assign addr[9745]= 2145835515;
assign addr[9746]= 2147470025;
assign addr[9747]= 2146380306;
assign addr[9748]= 2142567738;
assign addr[9749]= 2136037160;
assign addr[9750]= 2126796855;
assign addr[9751]= 2114858546;
assign addr[9752]= 2100237377;
assign addr[9753]= 2082951896;
assign addr[9754]= 2063024031;
assign addr[9755]= 2040479063;
assign addr[9756]= 2015345591;
assign addr[9757]= 1987655498;
assign addr[9758]= 1957443913;
assign addr[9759]= 1924749160;
assign addr[9760]= 1889612716;
assign addr[9761]= 1852079154;
assign addr[9762]= 1812196087;
assign addr[9763]= 1770014111;
assign addr[9764]= 1725586737;
assign addr[9765]= 1678970324;
assign addr[9766]= 1630224009;
assign addr[9767]= 1579409630;
assign addr[9768]= 1526591649;
assign addr[9769]= 1471837070;
assign addr[9770]= 1415215352;
assign addr[9771]= 1356798326;
assign addr[9772]= 1296660098;
assign addr[9773]= 1234876957;
assign addr[9774]= 1171527280;
assign addr[9775]= 1106691431;
assign addr[9776]= 1040451659;
assign addr[9777]= 972891995;
assign addr[9778]= 904098143;
assign addr[9779]= 834157373;
assign addr[9780]= 763158411;
assign addr[9781]= 691191324;
assign addr[9782]= 618347408;
assign addr[9783]= 544719071;
assign addr[9784]= 470399716;
assign addr[9785]= 395483624;
assign addr[9786]= 320065829;
assign addr[9787]= 244242007;
assign addr[9788]= 168108346;
assign addr[9789]= 91761426;
assign addr[9790]= 15298099;
assign addr[9791]= -61184634;
assign addr[9792]= -137589750;
assign addr[9793]= -213820322;
assign addr[9794]= -289779648;
assign addr[9795]= -365371365;
assign addr[9796]= -440499581;
assign addr[9797]= -515068990;
assign addr[9798]= -588984994;
assign addr[9799]= -662153826;
assign addr[9800]= -734482665;
assign addr[9801]= -805879757;
assign addr[9802]= -876254528;
assign addr[9803]= -945517704;
assign addr[9804]= -1013581418;
assign addr[9805]= -1080359326;
assign addr[9806]= -1145766716;
assign addr[9807]= -1209720613;
assign addr[9808]= -1272139887;
assign addr[9809]= -1332945355;
assign addr[9810]= -1392059879;
assign addr[9811]= -1449408469;
assign addr[9812]= -1504918373;
assign addr[9813]= -1558519173;
assign addr[9814]= -1610142873;
assign addr[9815]= -1659723983;
assign addr[9816]= -1707199606;
assign addr[9817]= -1752509516;
assign addr[9818]= -1795596234;
assign addr[9819]= -1836405100;
assign addr[9820]= -1874884346;
assign addr[9821]= -1910985158;
assign addr[9822]= -1944661739;
assign addr[9823]= -1975871368;
assign addr[9824]= -2004574453;
assign addr[9825]= -2030734582;
assign addr[9826]= -2054318569;
assign addr[9827]= -2075296495;
assign addr[9828]= -2093641749;
assign addr[9829]= -2109331059;
assign addr[9830]= -2122344521;
assign addr[9831]= -2132665626;
assign addr[9832]= -2140281282;
assign addr[9833]= -2145181827;
assign addr[9834]= -2147361045;
assign addr[9835]= -2146816171;
assign addr[9836]= -2143547897;
assign addr[9837]= -2137560369;
assign addr[9838]= -2128861181;
assign addr[9839]= -2117461370;
assign addr[9840]= -2103375398;
assign addr[9841]= -2086621133;
assign addr[9842]= -2067219829;
assign addr[9843]= -2045196100;
assign addr[9844]= -2020577882;
assign addr[9845]= -1993396407;
assign addr[9846]= -1963686155;
assign addr[9847]= -1931484818;
assign addr[9848]= -1896833245;
assign addr[9849]= -1859775393;
assign addr[9850]= -1820358275;
assign addr[9851]= -1778631892;
assign addr[9852]= -1734649179;
assign addr[9853]= -1688465931;
assign addr[9854]= -1640140734;
assign addr[9855]= -1589734894;
assign addr[9856]= -1537312353;
assign addr[9857]= -1482939614;
assign addr[9858]= -1426685652;
assign addr[9859]= -1368621831;
assign addr[9860]= -1308821808;
assign addr[9861]= -1247361445;
assign addr[9862]= -1184318708;
assign addr[9863]= -1119773573;
assign addr[9864]= -1053807919;
assign addr[9865]= -986505429;
assign addr[9866]= -917951481;
assign addr[9867]= -848233042;
assign addr[9868]= -777438554;
assign addr[9869]= -705657826;
assign addr[9870]= -632981917;
assign addr[9871]= -559503022;
assign addr[9872]= -485314355;
assign addr[9873]= -410510029;
assign addr[9874]= -335184940;
assign addr[9875]= -259434643;
assign addr[9876]= -183355234;
assign addr[9877]= -107043224;
assign addr[9878]= -30595422;
assign addr[9879]= 45891193;
assign addr[9880]= 122319591;
assign addr[9881]= 198592817;
assign addr[9882]= 274614114;
assign addr[9883]= 350287041;
assign addr[9884]= 425515602;
assign addr[9885]= 500204365;
assign addr[9886]= 574258580;
assign addr[9887]= 647584304;
assign addr[9888]= 720088517;
assign addr[9889]= 791679244;
assign addr[9890]= 862265664;
assign addr[9891]= 931758235;
assign addr[9892]= 1000068799;
assign addr[9893]= 1067110699;
assign addr[9894]= 1132798888;
assign addr[9895]= 1197050035;
assign addr[9896]= 1259782632;
assign addr[9897]= 1320917099;
assign addr[9898]= 1380375881;
assign addr[9899]= 1438083551;
assign addr[9900]= 1493966902;
assign addr[9901]= 1547955041;
assign addr[9902]= 1599979481;
assign addr[9903]= 1649974225;
assign addr[9904]= 1697875851;
assign addr[9905]= 1743623590;
assign addr[9906]= 1787159411;
assign addr[9907]= 1828428082;
assign addr[9908]= 1867377253;
assign addr[9909]= 1903957513;
assign addr[9910]= 1938122457;
assign addr[9911]= 1969828744;
assign addr[9912]= 1999036154;
assign addr[9913]= 2025707632;
assign addr[9914]= 2049809346;
assign addr[9915]= 2071310720;
assign addr[9916]= 2090184478;
assign addr[9917]= 2106406677;
assign addr[9918]= 2119956737;
assign addr[9919]= 2130817471;
assign addr[9920]= 2138975100;
assign addr[9921]= 2144419275;
assign addr[9922]= 2147143090;
assign addr[9923]= 2147143090;
assign addr[9924]= 2144419275;
assign addr[9925]= 2138975100;
assign addr[9926]= 2130817471;
assign addr[9927]= 2119956737;
assign addr[9928]= 2106406677;
assign addr[9929]= 2090184478;
assign addr[9930]= 2071310720;
assign addr[9931]= 2049809346;
assign addr[9932]= 2025707632;
assign addr[9933]= 1999036154;
assign addr[9934]= 1969828744;
assign addr[9935]= 1938122457;
assign addr[9936]= 1903957513;
assign addr[9937]= 1867377253;
assign addr[9938]= 1828428082;
assign addr[9939]= 1787159411;
assign addr[9940]= 1743623590;
assign addr[9941]= 1697875851;
assign addr[9942]= 1649974225;
assign addr[9943]= 1599979481;
assign addr[9944]= 1547955041;
assign addr[9945]= 1493966902;
assign addr[9946]= 1438083551;
assign addr[9947]= 1380375881;
assign addr[9948]= 1320917099;
assign addr[9949]= 1259782632;
assign addr[9950]= 1197050035;
assign addr[9951]= 1132798888;
assign addr[9952]= 1067110699;
assign addr[9953]= 1000068799;
assign addr[9954]= 931758235;
assign addr[9955]= 862265664;
assign addr[9956]= 791679244;
assign addr[9957]= 720088517;
assign addr[9958]= 647584304;
assign addr[9959]= 574258580;
assign addr[9960]= 500204365;
assign addr[9961]= 425515602;
assign addr[9962]= 350287041;
assign addr[9963]= 274614114;
assign addr[9964]= 198592817;
assign addr[9965]= 122319591;
assign addr[9966]= 45891193;
assign addr[9967]= -30595422;
assign addr[9968]= -107043224;
assign addr[9969]= -183355234;
assign addr[9970]= -259434643;
assign addr[9971]= -335184940;
assign addr[9972]= -410510029;
assign addr[9973]= -485314355;
assign addr[9974]= -559503022;
assign addr[9975]= -632981917;
assign addr[9976]= -705657826;
assign addr[9977]= -777438554;
assign addr[9978]= -848233042;
assign addr[9979]= -917951481;
assign addr[9980]= -986505429;
assign addr[9981]= -1053807919;
assign addr[9982]= -1119773573;
assign addr[9983]= -1184318708;
assign addr[9984]= -1247361445;
assign addr[9985]= -1308821808;
assign addr[9986]= -1368621831;
assign addr[9987]= -1426685652;
assign addr[9988]= -1482939614;
assign addr[9989]= -1537312353;
assign addr[9990]= -1589734894;
assign addr[9991]= -1640140734;
assign addr[9992]= -1688465931;
assign addr[9993]= -1734649179;
assign addr[9994]= -1778631892;
assign addr[9995]= -1820358275;
assign addr[9996]= -1859775393;
assign addr[9997]= -1896833245;
assign addr[9998]= -1931484818;
assign addr[9999]= -1963686155;
assign addr[10000]= -1993396407;
assign addr[10001]= -2020577882;
assign addr[10002]= -2045196100;
assign addr[10003]= -2067219829;
assign addr[10004]= -2086621133;
assign addr[10005]= -2103375398;
assign addr[10006]= -2117461370;
assign addr[10007]= -2128861181;
assign addr[10008]= -2137560369;
assign addr[10009]= -2143547897;
assign addr[10010]= -2146816171;
assign addr[10011]= -2147361045;
assign addr[10012]= -2145181827;
assign addr[10013]= -2140281282;
assign addr[10014]= -2132665626;
assign addr[10015]= -2122344521;
assign addr[10016]= -2109331059;
assign addr[10017]= -2093641749;
assign addr[10018]= -2075296495;
assign addr[10019]= -2054318569;
assign addr[10020]= -2030734582;
assign addr[10021]= -2004574453;
assign addr[10022]= -1975871368;
assign addr[10023]= -1944661739;
assign addr[10024]= -1910985158;
assign addr[10025]= -1874884346;
assign addr[10026]= -1836405100;
assign addr[10027]= -1795596234;
assign addr[10028]= -1752509516;
assign addr[10029]= -1707199606;
assign addr[10030]= -1659723983;
assign addr[10031]= -1610142873;
assign addr[10032]= -1558519173;
assign addr[10033]= -1504918373;
assign addr[10034]= -1449408469;
assign addr[10035]= -1392059879;
assign addr[10036]= -1332945355;
assign addr[10037]= -1272139887;
assign addr[10038]= -1209720613;
assign addr[10039]= -1145766716;
assign addr[10040]= -1080359326;
assign addr[10041]= -1013581418;
assign addr[10042]= -945517704;
assign addr[10043]= -876254528;
assign addr[10044]= -805879757;
assign addr[10045]= -734482665;
assign addr[10046]= -662153826;
assign addr[10047]= -588984994;
assign addr[10048]= -515068990;
assign addr[10049]= -440499581;
assign addr[10050]= -365371365;
assign addr[10051]= -289779648;
assign addr[10052]= -213820322;
assign addr[10053]= -137589750;
assign addr[10054]= -61184634;
assign addr[10055]= 15298099;
assign addr[10056]= 91761426;
assign addr[10057]= 168108346;
assign addr[10058]= 244242007;
assign addr[10059]= 320065829;
assign addr[10060]= 395483624;
assign addr[10061]= 470399716;
assign addr[10062]= 544719071;
assign addr[10063]= 618347408;
assign addr[10064]= 691191324;
assign addr[10065]= 763158411;
assign addr[10066]= 834157373;
assign addr[10067]= 904098143;
assign addr[10068]= 972891995;
assign addr[10069]= 1040451659;
assign addr[10070]= 1106691431;
assign addr[10071]= 1171527280;
assign addr[10072]= 1234876957;
assign addr[10073]= 1296660098;
assign addr[10074]= 1356798326;
assign addr[10075]= 1415215352;
assign addr[10076]= 1471837070;
assign addr[10077]= 1526591649;
assign addr[10078]= 1579409630;
assign addr[10079]= 1630224009;
assign addr[10080]= 1678970324;
assign addr[10081]= 1725586737;
assign addr[10082]= 1770014111;
assign addr[10083]= 1812196087;
assign addr[10084]= 1852079154;
assign addr[10085]= 1889612716;
assign addr[10086]= 1924749160;
assign addr[10087]= 1957443913;
assign addr[10088]= 1987655498;
assign addr[10089]= 2015345591;
assign addr[10090]= 2040479063;
assign addr[10091]= 2063024031;
assign addr[10092]= 2082951896;
assign addr[10093]= 2100237377;
assign addr[10094]= 2114858546;
assign addr[10095]= 2126796855;
assign addr[10096]= 2136037160;
assign addr[10097]= 2142567738;
assign addr[10098]= 2146380306;
assign addr[10099]= 2147470025;
assign addr[10100]= 2145835515;
assign addr[10101]= 2141478848;
assign addr[10102]= 2134405552;
assign addr[10103]= 2124624598;
assign addr[10104]= 2112148396;
assign addr[10105]= 2096992772;
assign addr[10106]= 2079176953;
assign addr[10107]= 2058723538;
assign addr[10108]= 2035658475;
assign addr[10109]= 2010011024;
assign addr[10110]= 1981813720;
assign addr[10111]= 1951102334;
assign addr[10112]= 1917915825;
assign addr[10113]= 1882296293;
assign addr[10114]= 1844288924;
assign addr[10115]= 1803941934;
assign addr[10116]= 1761306505;
assign addr[10117]= 1716436725;
assign addr[10118]= 1669389513;
assign addr[10119]= 1620224553;
assign addr[10120]= 1569004214;
assign addr[10121]= 1515793473;
assign addr[10122]= 1460659832;
assign addr[10123]= 1403673233;
assign addr[10124]= 1344905966;
assign addr[10125]= 1284432584;
assign addr[10126]= 1222329801;
assign addr[10127]= 1158676398;
assign addr[10128]= 1093553126;
assign addr[10129]= 1027042599;
assign addr[10130]= 959229189;
assign addr[10131]= 890198924;
assign addr[10132]= 820039373;
assign addr[10133]= 748839539;
assign addr[10134]= 676689746;
assign addr[10135]= 603681519;
assign addr[10136]= 529907477;
assign addr[10137]= 455461206;
assign addr[10138]= 380437148;
assign addr[10139]= 304930476;
assign addr[10140]= 229036977;
assign addr[10141]= 152852926;
assign addr[10142]= 76474970;
assign addr[10143]= 0;
assign addr[10144]= -76474970;
assign addr[10145]= -152852926;
assign addr[10146]= -229036977;
assign addr[10147]= -304930476;
assign addr[10148]= -380437148;
assign addr[10149]= -455461206;
assign addr[10150]= -529907477;
assign addr[10151]= -603681519;
assign addr[10152]= -676689746;
assign addr[10153]= -748839539;
assign addr[10154]= -820039373;
assign addr[10155]= -890198924;
assign addr[10156]= -959229189;
assign addr[10157]= -1027042599;
assign addr[10158]= -1093553126;
assign addr[10159]= -1158676398;
assign addr[10160]= -1222329801;
assign addr[10161]= -1284432584;
assign addr[10162]= -1344905966;
assign addr[10163]= -1403673233;
assign addr[10164]= -1460659832;
assign addr[10165]= -1515793473;
assign addr[10166]= -1569004214;
assign addr[10167]= -1620224553;
assign addr[10168]= -1669389513;
assign addr[10169]= -1716436725;
assign addr[10170]= -1761306505;
assign addr[10171]= -1803941934;
assign addr[10172]= -1844288924;
assign addr[10173]= -1882296293;
assign addr[10174]= -1917915825;
assign addr[10175]= -1951102334;
assign addr[10176]= -1981813720;
assign addr[10177]= -2010011024;
assign addr[10178]= -2035658475;
assign addr[10179]= -2058723538;
assign addr[10180]= -2079176953;
assign addr[10181]= -2096992772;
assign addr[10182]= -2112148396;
assign addr[10183]= -2124624598;
assign addr[10184]= -2134405552;
assign addr[10185]= -2141478848;
assign addr[10186]= -2145835515;
assign addr[10187]= -2147470025;
assign addr[10188]= -2146380306;
assign addr[10189]= -2142567738;
assign addr[10190]= -2136037160;
assign addr[10191]= -2126796855;
assign addr[10192]= -2114858546;
assign addr[10193]= -2100237377;
assign addr[10194]= -2082951896;
assign addr[10195]= -2063024031;
assign addr[10196]= -2040479063;
assign addr[10197]= -2015345591;
assign addr[10198]= -1987655498;
assign addr[10199]= -1957443913;
assign addr[10200]= -1924749160;
assign addr[10201]= -1889612716;
assign addr[10202]= -1852079154;
assign addr[10203]= -1812196087;
assign addr[10204]= -1770014111;
assign addr[10205]= -1725586737;
assign addr[10206]= -1678970324;
assign addr[10207]= -1630224009;
assign addr[10208]= -1579409630;
assign addr[10209]= -1526591649;
assign addr[10210]= -1471837070;
assign addr[10211]= -1415215352;
assign addr[10212]= -1356798326;
assign addr[10213]= -1296660098;
assign addr[10214]= -1234876957;
assign addr[10215]= -1171527280;
assign addr[10216]= -1106691431;
assign addr[10217]= -1040451659;
assign addr[10218]= -972891995;
assign addr[10219]= -904098143;
assign addr[10220]= -834157373;
assign addr[10221]= -763158411;
assign addr[10222]= -691191324;
assign addr[10223]= -618347408;
assign addr[10224]= -544719071;
assign addr[10225]= -470399716;
assign addr[10226]= -395483624;
assign addr[10227]= -320065829;
assign addr[10228]= -244242007;
assign addr[10229]= -168108346;
assign addr[10230]= -91761426;
assign addr[10231]= -15298099;
assign addr[10232]= 61184634;
assign addr[10233]= 137589750;
assign addr[10234]= 213820322;
assign addr[10235]= 289779648;
assign addr[10236]= 365371365;
assign addr[10237]= 440499581;
assign addr[10238]= 515068990;
assign addr[10239]= 588984994;
assign addr[10240]= 662153826;
assign addr[10241]= 734482665;
assign addr[10242]= 805879757;
assign addr[10243]= 876254528;
assign addr[10244]= 945517704;
assign addr[10245]= 1013581418;
assign addr[10246]= 1080359326;
assign addr[10247]= 1145766716;
assign addr[10248]= 1209720613;
assign addr[10249]= 1272139887;
assign addr[10250]= 1332945355;
assign addr[10251]= 1392059879;
assign addr[10252]= 1449408469;
assign addr[10253]= 1504918373;
assign addr[10254]= 1558519173;
assign addr[10255]= 1610142873;
assign addr[10256]= 1659723983;
assign addr[10257]= 1707199606;
assign addr[10258]= 1752509516;
assign addr[10259]= 1795596234;
assign addr[10260]= 1836405100;
assign addr[10261]= 1874884346;
assign addr[10262]= 1910985158;
assign addr[10263]= 1944661739;
assign addr[10264]= 1975871368;
assign addr[10265]= 2004574453;
assign addr[10266]= 2030734582;
assign addr[10267]= 2054318569;
assign addr[10268]= 2075296495;
assign addr[10269]= 2093641749;
assign addr[10270]= 2109331059;
assign addr[10271]= 2122344521;
assign addr[10272]= 2132665626;
assign addr[10273]= 2140281282;
assign addr[10274]= 2145181827;
assign addr[10275]= 2147361045;
assign addr[10276]= 2146816171;
assign addr[10277]= 2143547897;
assign addr[10278]= 2137560369;
assign addr[10279]= 2128861181;
assign addr[10280]= 2117461370;
assign addr[10281]= 2103375398;
assign addr[10282]= 2086621133;
assign addr[10283]= 2067219829;
assign addr[10284]= 2045196100;
assign addr[10285]= 2020577882;
assign addr[10286]= 1993396407;
assign addr[10287]= 1963686155;
assign addr[10288]= 1931484818;
assign addr[10289]= 1896833245;
assign addr[10290]= 1859775393;
assign addr[10291]= 1820358275;
assign addr[10292]= 1778631892;
assign addr[10293]= 1734649179;
assign addr[10294]= 1688465931;
assign addr[10295]= 1640140734;
assign addr[10296]= 1589734894;
assign addr[10297]= 1537312353;
assign addr[10298]= 1482939614;
assign addr[10299]= 1426685652;
assign addr[10300]= 1368621831;
assign addr[10301]= 1308821808;
assign addr[10302]= 1247361445;
assign addr[10303]= 1184318708;
assign addr[10304]= 1119773573;
assign addr[10305]= 1053807919;
assign addr[10306]= 986505429;
assign addr[10307]= 917951481;
assign addr[10308]= 848233042;
assign addr[10309]= 777438554;
assign addr[10310]= 705657826;
assign addr[10311]= 632981917;
assign addr[10312]= 559503022;
assign addr[10313]= 485314355;
assign addr[10314]= 410510029;
assign addr[10315]= 335184940;
assign addr[10316]= 259434643;
assign addr[10317]= 183355234;
assign addr[10318]= 107043224;
assign addr[10319]= 30595422;
assign addr[10320]= -45891193;
assign addr[10321]= -122319591;
assign addr[10322]= -198592817;
assign addr[10323]= -274614114;
assign addr[10324]= -350287041;
assign addr[10325]= -425515602;
assign addr[10326]= -500204365;
assign addr[10327]= -574258580;
assign addr[10328]= -647584304;
assign addr[10329]= -720088517;
assign addr[10330]= -791679244;
assign addr[10331]= -862265664;
assign addr[10332]= -931758235;
assign addr[10333]= -1000068799;
assign addr[10334]= -1067110699;
assign addr[10335]= -1132798888;
assign addr[10336]= -1197050035;
assign addr[10337]= -1259782632;
assign addr[10338]= -1320917099;
assign addr[10339]= -1380375881;
assign addr[10340]= -1438083551;
assign addr[10341]= -1493966902;
assign addr[10342]= -1547955041;
assign addr[10343]= -1599979481;
assign addr[10344]= -1649974225;
assign addr[10345]= -1697875851;
assign addr[10346]= -1743623590;
assign addr[10347]= -1787159411;
assign addr[10348]= -1828428082;
assign addr[10349]= -1867377253;
assign addr[10350]= -1903957513;
assign addr[10351]= -1938122457;
assign addr[10352]= -1969828744;
assign addr[10353]= -1999036154;
assign addr[10354]= -2025707632;
assign addr[10355]= -2049809346;
assign addr[10356]= -2071310720;
assign addr[10357]= -2090184478;
assign addr[10358]= -2106406677;
assign addr[10359]= -2119956737;
assign addr[10360]= -2130817471;
assign addr[10361]= -2138975100;
assign addr[10362]= -2144419275;
assign addr[10363]= -2147143090;
assign addr[10364]= -2147143090;
assign addr[10365]= -2144419275;
assign addr[10366]= -2138975100;
assign addr[10367]= -2130817471;
assign addr[10368]= -2119956737;
assign addr[10369]= -2106406677;
assign addr[10370]= -2090184478;
assign addr[10371]= -2071310720;
assign addr[10372]= -2049809346;
assign addr[10373]= -2025707632;
assign addr[10374]= -1999036154;
assign addr[10375]= -1969828744;
assign addr[10376]= -1938122457;
assign addr[10377]= -1903957513;
assign addr[10378]= -1867377253;
assign addr[10379]= -1828428082;
assign addr[10380]= -1787159411;
assign addr[10381]= -1743623590;
assign addr[10382]= -1697875851;
assign addr[10383]= -1649974225;
assign addr[10384]= -1599979481;
assign addr[10385]= -1547955041;
assign addr[10386]= -1493966902;
assign addr[10387]= -1438083551;
assign addr[10388]= -1380375881;
assign addr[10389]= -1320917099;
assign addr[10390]= -1259782632;
assign addr[10391]= -1197050035;
assign addr[10392]= -1132798888;
assign addr[10393]= -1067110699;
assign addr[10394]= -1000068799;
assign addr[10395]= -931758235;
assign addr[10396]= -862265664;
assign addr[10397]= -791679244;
assign addr[10398]= -720088517;
assign addr[10399]= -647584304;
assign addr[10400]= -574258580;
assign addr[10401]= -500204365;
assign addr[10402]= -425515602;
assign addr[10403]= -350287041;
assign addr[10404]= -274614114;
assign addr[10405]= -198592817;
assign addr[10406]= -122319591;
assign addr[10407]= -45891193;
assign addr[10408]= 30595422;
assign addr[10409]= 107043224;
assign addr[10410]= 183355234;
assign addr[10411]= 259434643;
assign addr[10412]= 335184940;
assign addr[10413]= 410510029;
assign addr[10414]= 485314355;
assign addr[10415]= 559503022;
assign addr[10416]= 632981917;
assign addr[10417]= 705657826;
assign addr[10418]= 777438554;
assign addr[10419]= 848233042;
assign addr[10420]= 917951481;
assign addr[10421]= 986505429;
assign addr[10422]= 1053807919;
assign addr[10423]= 1119773573;
assign addr[10424]= 1184318708;
assign addr[10425]= 1247361445;
assign addr[10426]= 1308821808;
assign addr[10427]= 1368621831;
assign addr[10428]= 1426685652;
assign addr[10429]= 1482939614;
assign addr[10430]= 1537312353;
assign addr[10431]= 1589734894;
assign addr[10432]= 1640140734;
assign addr[10433]= 1688465931;
assign addr[10434]= 1734649179;
assign addr[10435]= 1778631892;
assign addr[10436]= 1820358275;
assign addr[10437]= 1859775393;
assign addr[10438]= 1896833245;
assign addr[10439]= 1931484818;
assign addr[10440]= 1963686155;
assign addr[10441]= 1993396407;
assign addr[10442]= 2020577882;
assign addr[10443]= 2045196100;
assign addr[10444]= 2067219829;
assign addr[10445]= 2086621133;
assign addr[10446]= 2103375398;
assign addr[10447]= 2117461370;
assign addr[10448]= 2128861181;
assign addr[10449]= 2137560369;
assign addr[10450]= 2143547897;
assign addr[10451]= 2146816171;
assign addr[10452]= 2147361045;
assign addr[10453]= 2145181827;
assign addr[10454]= 2140281282;
assign addr[10455]= 2132665626;
assign addr[10456]= 2122344521;
assign addr[10457]= 2109331059;
assign addr[10458]= 2093641749;
assign addr[10459]= 2075296495;
assign addr[10460]= 2054318569;
assign addr[10461]= 2030734582;
assign addr[10462]= 2004574453;
assign addr[10463]= 1975871368;
assign addr[10464]= 1944661739;
assign addr[10465]= 1910985158;
assign addr[10466]= 1874884346;
assign addr[10467]= 1836405100;
assign addr[10468]= 1795596234;
assign addr[10469]= 1752509516;
assign addr[10470]= 1707199606;
assign addr[10471]= 1659723983;
assign addr[10472]= 1610142873;
assign addr[10473]= 1558519173;
assign addr[10474]= 1504918373;
assign addr[10475]= 1449408469;
assign addr[10476]= 1392059879;
assign addr[10477]= 1332945355;
assign addr[10478]= 1272139887;
assign addr[10479]= 1209720613;
assign addr[10480]= 1145766716;
assign addr[10481]= 1080359326;
assign addr[10482]= 1013581418;
assign addr[10483]= 945517704;
assign addr[10484]= 876254528;
assign addr[10485]= 805879757;
assign addr[10486]= 734482665;
assign addr[10487]= 662153826;
assign addr[10488]= 588984994;
assign addr[10489]= 515068990;
assign addr[10490]= 440499581;
assign addr[10491]= 365371365;
assign addr[10492]= 289779648;
assign addr[10493]= 213820322;
assign addr[10494]= 137589750;
assign addr[10495]= 61184634;
assign addr[10496]= -15298099;
assign addr[10497]= -91761426;
assign addr[10498]= -168108346;
assign addr[10499]= -244242007;
assign addr[10500]= -320065829;
assign addr[10501]= -395483624;
assign addr[10502]= -470399716;
assign addr[10503]= -544719071;
assign addr[10504]= -618347408;
assign addr[10505]= -691191324;
assign addr[10506]= -763158411;
assign addr[10507]= -834157373;
assign addr[10508]= -904098143;
assign addr[10509]= -972891995;
assign addr[10510]= -1040451659;
assign addr[10511]= -1106691431;
assign addr[10512]= -1171527280;
assign addr[10513]= -1234876957;
assign addr[10514]= -1296660098;
assign addr[10515]= -1356798326;
assign addr[10516]= -1415215352;
assign addr[10517]= -1471837070;
assign addr[10518]= -1526591649;
assign addr[10519]= -1579409630;
assign addr[10520]= -1630224009;
assign addr[10521]= -1678970324;
assign addr[10522]= -1725586737;
assign addr[10523]= -1770014111;
assign addr[10524]= -1812196087;
assign addr[10525]= -1852079154;
assign addr[10526]= -1889612716;
assign addr[10527]= -1924749160;
assign addr[10528]= -1957443913;
assign addr[10529]= -1987655498;
assign addr[10530]= -2015345591;
assign addr[10531]= -2040479063;
assign addr[10532]= -2063024031;
assign addr[10533]= -2082951896;
assign addr[10534]= -2100237377;
assign addr[10535]= -2114858546;
assign addr[10536]= -2126796855;
assign addr[10537]= -2136037160;
assign addr[10538]= -2142567738;
assign addr[10539]= -2146380306;
assign addr[10540]= -2147470025;
assign addr[10541]= -2145835515;
assign addr[10542]= -2141478848;
assign addr[10543]= -2134405552;
assign addr[10544]= -2124624598;
assign addr[10545]= -2112148396;
assign addr[10546]= -2096992772;
assign addr[10547]= -2079176953;
assign addr[10548]= -2058723538;
assign addr[10549]= -2035658475;
assign addr[10550]= -2010011024;
assign addr[10551]= -1981813720;
assign addr[10552]= -1951102334;
assign addr[10553]= -1917915825;
assign addr[10554]= -1882296293;
assign addr[10555]= -1844288924;
assign addr[10556]= -1803941934;
assign addr[10557]= -1761306505;
assign addr[10558]= -1716436725;
assign addr[10559]= -1669389513;
assign addr[10560]= -1620224553;
assign addr[10561]= -1569004214;
assign addr[10562]= -1515793473;
assign addr[10563]= -1460659832;
assign addr[10564]= -1403673233;
assign addr[10565]= -1344905966;
assign addr[10566]= -1284432584;
assign addr[10567]= -1222329801;
assign addr[10568]= -1158676398;
assign addr[10569]= -1093553126;
assign addr[10570]= -1027042599;
assign addr[10571]= -959229189;
assign addr[10572]= -890198924;
assign addr[10573]= -820039373;
assign addr[10574]= -748839539;
assign addr[10575]= -676689746;
assign addr[10576]= -603681519;
assign addr[10577]= -529907477;
assign addr[10578]= -455461206;
assign addr[10579]= -380437148;
assign addr[10580]= -304930476;
assign addr[10581]= -229036977;
assign addr[10582]= -152852926;
assign addr[10583]= -76474970;
assign addr[10584]= 0;
assign addr[10585]= 76474970;
assign addr[10586]= 152852926;
assign addr[10587]= 229036977;
assign addr[10588]= 304930476;
assign addr[10589]= 380437148;
assign addr[10590]= 455461206;
assign addr[10591]= 529907477;
assign addr[10592]= 603681519;
assign addr[10593]= 676689746;
assign addr[10594]= 748839539;
assign addr[10595]= 820039373;
assign addr[10596]= 890198924;
assign addr[10597]= 959229189;
assign addr[10598]= 1027042599;
assign addr[10599]= 1093553126;
assign addr[10600]= 1158676398;
assign addr[10601]= 1222329801;
assign addr[10602]= 1284432584;
assign addr[10603]= 1344905966;
assign addr[10604]= 1403673233;
assign addr[10605]= 1460659832;
assign addr[10606]= 1515793473;
assign addr[10607]= 1569004214;
assign addr[10608]= 1620224553;
assign addr[10609]= 1669389513;
assign addr[10610]= 1716436725;
assign addr[10611]= 1761306505;
assign addr[10612]= 1803941934;
assign addr[10613]= 1844288924;
assign addr[10614]= 1882296293;
assign addr[10615]= 1917915825;
assign addr[10616]= 1951102334;
assign addr[10617]= 1981813720;
assign addr[10618]= 2010011024;
assign addr[10619]= 2035658475;
assign addr[10620]= 2058723538;
assign addr[10621]= 2079176953;
assign addr[10622]= 2096992772;
assign addr[10623]= 2112148396;
assign addr[10624]= 2124624598;
assign addr[10625]= 2134405552;
assign addr[10626]= 2141478848;
assign addr[10627]= 2145835515;
assign addr[10628]= 2147470025;
assign addr[10629]= 2146380306;
assign addr[10630]= 2142567738;
assign addr[10631]= 2136037160;
assign addr[10632]= 2126796855;
assign addr[10633]= 2114858546;
assign addr[10634]= 2100237377;
assign addr[10635]= 2082951896;
assign addr[10636]= 2063024031;
assign addr[10637]= 2040479063;
assign addr[10638]= 2015345591;
assign addr[10639]= 1987655498;
assign addr[10640]= 1957443913;
assign addr[10641]= 1924749160;
assign addr[10642]= 1889612716;
assign addr[10643]= 1852079154;
assign addr[10644]= 1812196087;
assign addr[10645]= 1770014111;
assign addr[10646]= 1725586737;
assign addr[10647]= 1678970324;
assign addr[10648]= 1630224009;
assign addr[10649]= 1579409630;
assign addr[10650]= 1526591649;
assign addr[10651]= 1471837070;
assign addr[10652]= 1415215352;
assign addr[10653]= 1356798326;
assign addr[10654]= 1296660098;
assign addr[10655]= 1234876957;
assign addr[10656]= 1171527280;
assign addr[10657]= 1106691431;
assign addr[10658]= 1040451659;
assign addr[10659]= 972891995;
assign addr[10660]= 904098143;
assign addr[10661]= 834157373;
assign addr[10662]= 763158411;
assign addr[10663]= 691191324;
assign addr[10664]= 618347408;
assign addr[10665]= 544719071;
assign addr[10666]= 470399716;
assign addr[10667]= 395483624;
assign addr[10668]= 320065829;
assign addr[10669]= 244242007;
assign addr[10670]= 168108346;
assign addr[10671]= 91761426;
assign addr[10672]= 15298099;
assign addr[10673]= -61184634;
assign addr[10674]= -137589750;
assign addr[10675]= -213820322;
assign addr[10676]= -289779648;
assign addr[10677]= -365371365;
assign addr[10678]= -440499581;
assign addr[10679]= -515068990;
assign addr[10680]= -588984994;
assign addr[10681]= -662153826;
assign addr[10682]= -734482665;
assign addr[10683]= -805879757;
assign addr[10684]= -876254528;
assign addr[10685]= -945517704;
assign addr[10686]= -1013581418;
assign addr[10687]= -1080359326;
assign addr[10688]= -1145766716;
assign addr[10689]= -1209720613;
assign addr[10690]= -1272139887;
assign addr[10691]= -1332945355;
assign addr[10692]= -1392059879;
assign addr[10693]= -1449408469;
assign addr[10694]= -1504918373;
assign addr[10695]= -1558519173;
assign addr[10696]= -1610142873;
assign addr[10697]= -1659723983;
assign addr[10698]= -1707199606;
assign addr[10699]= -1752509516;
assign addr[10700]= -1795596234;
assign addr[10701]= -1836405100;
assign addr[10702]= -1874884346;
assign addr[10703]= -1910985158;
assign addr[10704]= -1944661739;
assign addr[10705]= -1975871368;
assign addr[10706]= -2004574453;
assign addr[10707]= -2030734582;
assign addr[10708]= -2054318569;
assign addr[10709]= -2075296495;
assign addr[10710]= -2093641749;
assign addr[10711]= -2109331059;
assign addr[10712]= -2122344521;
assign addr[10713]= -2132665626;
assign addr[10714]= -2140281282;
assign addr[10715]= -2145181827;
assign addr[10716]= -2147361045;
assign addr[10717]= -2146816171;
assign addr[10718]= -2143547897;
assign addr[10719]= -2137560369;
assign addr[10720]= -2128861181;
assign addr[10721]= -2117461370;
assign addr[10722]= -2103375398;
assign addr[10723]= -2086621133;
assign addr[10724]= -2067219829;
assign addr[10725]= -2045196100;
assign addr[10726]= -2020577882;
assign addr[10727]= -1993396407;
assign addr[10728]= -1963686155;
assign addr[10729]= -1931484818;
assign addr[10730]= -1896833245;
assign addr[10731]= -1859775393;
assign addr[10732]= -1820358275;
assign addr[10733]= -1778631892;
assign addr[10734]= -1734649179;
assign addr[10735]= -1688465931;
assign addr[10736]= -1640140734;
assign addr[10737]= -1589734894;
assign addr[10738]= -1537312353;
assign addr[10739]= -1482939614;
assign addr[10740]= -1426685652;
assign addr[10741]= -1368621831;
assign addr[10742]= -1308821808;
assign addr[10743]= -1247361445;
assign addr[10744]= -1184318708;
assign addr[10745]= -1119773573;
assign addr[10746]= -1053807919;
assign addr[10747]= -986505429;
assign addr[10748]= -917951481;
assign addr[10749]= -848233042;
assign addr[10750]= -777438554;
assign addr[10751]= -705657826;
assign addr[10752]= -632981917;
assign addr[10753]= -559503022;
assign addr[10754]= -485314355;
assign addr[10755]= -410510029;
assign addr[10756]= -335184940;
assign addr[10757]= -259434643;
assign addr[10758]= -183355234;
assign addr[10759]= -107043224;
assign addr[10760]= -30595422;
assign addr[10761]= 45891193;
assign addr[10762]= 122319591;
assign addr[10763]= 198592817;
assign addr[10764]= 274614114;
assign addr[10765]= 350287041;
assign addr[10766]= 425515602;
assign addr[10767]= 500204365;
assign addr[10768]= 574258580;
assign addr[10769]= 647584304;
assign addr[10770]= 720088517;
assign addr[10771]= 791679244;
assign addr[10772]= 862265664;
assign addr[10773]= 931758235;
assign addr[10774]= 1000068799;
assign addr[10775]= 1067110699;
assign addr[10776]= 1132798888;
assign addr[10777]= 1197050035;
assign addr[10778]= 1259782632;
assign addr[10779]= 1320917099;
assign addr[10780]= 1380375881;
assign addr[10781]= 1438083551;
assign addr[10782]= 1493966902;
assign addr[10783]= 1547955041;
assign addr[10784]= 1599979481;
assign addr[10785]= 1649974225;
assign addr[10786]= 1697875851;
assign addr[10787]= 1743623590;
assign addr[10788]= 1787159411;
assign addr[10789]= 1828428082;
assign addr[10790]= 1867377253;
assign addr[10791]= 1903957513;
assign addr[10792]= 1938122457;
assign addr[10793]= 1969828744;
assign addr[10794]= 1999036154;
assign addr[10795]= 2025707632;
assign addr[10796]= 2049809346;
assign addr[10797]= 2071310720;
assign addr[10798]= 2090184478;
assign addr[10799]= 2106406677;
assign addr[10800]= 2119956737;
assign addr[10801]= 2130817471;
assign addr[10802]= 2138975100;
assign addr[10803]= 2144419275;
assign addr[10804]= 2147143090;
assign addr[10805]= 2147143090;
assign addr[10806]= 2144419275;
assign addr[10807]= 2138975100;
assign addr[10808]= 2130817471;
assign addr[10809]= 2119956737;
assign addr[10810]= 2106406677;
assign addr[10811]= 2090184478;
assign addr[10812]= 2071310720;
assign addr[10813]= 2049809346;
assign addr[10814]= 2025707632;
assign addr[10815]= 1999036154;
assign addr[10816]= 1969828744;
assign addr[10817]= 1938122457;
assign addr[10818]= 1903957513;
assign addr[10819]= 1867377253;
assign addr[10820]= 1828428082;
assign addr[10821]= 1787159411;
assign addr[10822]= 1743623590;
assign addr[10823]= 1697875851;
assign addr[10824]= 1649974225;
assign addr[10825]= 1599979481;
assign addr[10826]= 1547955041;
assign addr[10827]= 1493966902;
assign addr[10828]= 1438083551;
assign addr[10829]= 1380375881;
assign addr[10830]= 1320917099;
assign addr[10831]= 1259782632;
assign addr[10832]= 1197050035;
assign addr[10833]= 1132798888;
assign addr[10834]= 1067110699;
assign addr[10835]= 1000068799;
assign addr[10836]= 931758235;
assign addr[10837]= 862265664;
assign addr[10838]= 791679244;
assign addr[10839]= 720088517;
assign addr[10840]= 647584304;
assign addr[10841]= 574258580;
assign addr[10842]= 500204365;
assign addr[10843]= 425515602;
assign addr[10844]= 350287041;
assign addr[10845]= 274614114;
assign addr[10846]= 198592817;
assign addr[10847]= 122319591;
assign addr[10848]= 45891193;
assign addr[10849]= -30595422;
assign addr[10850]= -107043224;
assign addr[10851]= -183355234;
assign addr[10852]= -259434643;
assign addr[10853]= -335184940;
assign addr[10854]= -410510029;
assign addr[10855]= -485314355;
assign addr[10856]= -559503022;
assign addr[10857]= -632981917;
assign addr[10858]= -705657826;
assign addr[10859]= -777438554;
assign addr[10860]= -848233042;
assign addr[10861]= -917951481;
assign addr[10862]= -986505429;
assign addr[10863]= -1053807919;
assign addr[10864]= -1119773573;
assign addr[10865]= -1184318708;
assign addr[10866]= -1247361445;
assign addr[10867]= -1308821808;
assign addr[10868]= -1368621831;
assign addr[10869]= -1426685652;
assign addr[10870]= -1482939614;
assign addr[10871]= -1537312353;
assign addr[10872]= -1589734894;
assign addr[10873]= -1640140734;
assign addr[10874]= -1688465931;
assign addr[10875]= -1734649179;
assign addr[10876]= -1778631892;
assign addr[10877]= -1820358275;
assign addr[10878]= -1859775393;
assign addr[10879]= -1896833245;
assign addr[10880]= -1931484818;
assign addr[10881]= -1963686155;
assign addr[10882]= -1993396407;
assign addr[10883]= -2020577882;
assign addr[10884]= -2045196100;
assign addr[10885]= -2067219829;
assign addr[10886]= -2086621133;
assign addr[10887]= -2103375398;
assign addr[10888]= -2117461370;
assign addr[10889]= -2128861181;
assign addr[10890]= -2137560369;
assign addr[10891]= -2143547897;
assign addr[10892]= -2146816171;
assign addr[10893]= -2147361045;
assign addr[10894]= -2145181827;
assign addr[10895]= -2140281282;
assign addr[10896]= -2132665626;
assign addr[10897]= -2122344521;
assign addr[10898]= -2109331059;
assign addr[10899]= -2093641749;
assign addr[10900]= -2075296495;
assign addr[10901]= -2054318569;
assign addr[10902]= -2030734582;
assign addr[10903]= -2004574453;
assign addr[10904]= -1975871368;
assign addr[10905]= -1944661739;
assign addr[10906]= -1910985158;
assign addr[10907]= -1874884346;
assign addr[10908]= -1836405100;
assign addr[10909]= -1795596234;
assign addr[10910]= -1752509516;
assign addr[10911]= -1707199606;
assign addr[10912]= -1659723983;
assign addr[10913]= -1610142873;
assign addr[10914]= -1558519173;
assign addr[10915]= -1504918373;
assign addr[10916]= -1449408469;
assign addr[10917]= -1392059879;
assign addr[10918]= -1332945355;
assign addr[10919]= -1272139887;
assign addr[10920]= -1209720613;
assign addr[10921]= -1145766716;
assign addr[10922]= -1080359326;
assign addr[10923]= -1013581418;
assign addr[10924]= -945517704;
assign addr[10925]= -876254528;
assign addr[10926]= -805879757;
assign addr[10927]= -734482665;
assign addr[10928]= -662153826;
assign addr[10929]= -588984994;
assign addr[10930]= -515068990;
assign addr[10931]= -440499581;
assign addr[10932]= -365371365;
assign addr[10933]= -289779648;
assign addr[10934]= -213820322;
assign addr[10935]= -137589750;
assign addr[10936]= -61184634;
assign addr[10937]= 15298099;
assign addr[10938]= 91761426;
assign addr[10939]= 168108346;
assign addr[10940]= 244242007;
assign addr[10941]= 320065829;
assign addr[10942]= 395483624;
assign addr[10943]= 470399716;
assign addr[10944]= 544719071;
assign addr[10945]= 618347408;
assign addr[10946]= 691191324;
assign addr[10947]= 763158411;
assign addr[10948]= 834157373;
assign addr[10949]= 904098143;
assign addr[10950]= 972891995;
assign addr[10951]= 1040451659;
assign addr[10952]= 1106691431;
assign addr[10953]= 1171527280;
assign addr[10954]= 1234876957;
assign addr[10955]= 1296660098;
assign addr[10956]= 1356798326;
assign addr[10957]= 1415215352;
assign addr[10958]= 1471837070;
assign addr[10959]= 1526591649;
assign addr[10960]= 1579409630;
assign addr[10961]= 1630224009;
assign addr[10962]= 1678970324;
assign addr[10963]= 1725586737;
assign addr[10964]= 1770014111;
assign addr[10965]= 1812196087;
assign addr[10966]= 1852079154;
assign addr[10967]= 1889612716;
assign addr[10968]= 1924749160;
assign addr[10969]= 1957443913;
assign addr[10970]= 1987655498;
assign addr[10971]= 2015345591;
assign addr[10972]= 2040479063;
assign addr[10973]= 2063024031;
assign addr[10974]= 2082951896;
assign addr[10975]= 2100237377;
assign addr[10976]= 2114858546;
assign addr[10977]= 2126796855;
assign addr[10978]= 2136037160;
assign addr[10979]= 2142567738;
assign addr[10980]= 2146380306;
assign addr[10981]= 2147470025;
assign addr[10982]= 2145835515;
assign addr[10983]= 2141478848;
assign addr[10984]= 2134405552;
assign addr[10985]= 2124624598;
assign addr[10986]= 2112148396;
assign addr[10987]= 2096992772;
assign addr[10988]= 2079176953;
assign addr[10989]= 2058723538;
assign addr[10990]= 2035658475;
assign addr[10991]= 2010011024;
assign addr[10992]= 1981813720;
assign addr[10993]= 1951102334;
assign addr[10994]= 1917915825;
assign addr[10995]= 1882296293;
assign addr[10996]= 1844288924;
assign addr[10997]= 1803941934;
assign addr[10998]= 1761306505;
assign addr[10999]= 1716436725;
assign addr[11000]= 1669389513;
assign addr[11001]= 1620224553;
assign addr[11002]= 1569004214;
assign addr[11003]= 1515793473;
assign addr[11004]= 1460659832;
assign addr[11005]= 1403673233;
assign addr[11006]= 1344905966;
assign addr[11007]= 1284432584;
assign addr[11008]= 1222329801;
assign addr[11009]= 1158676398;
assign addr[11010]= 1093553126;
assign addr[11011]= 1027042599;
assign addr[11012]= 959229189;
assign addr[11013]= 890198924;
assign addr[11014]= 820039373;
assign addr[11015]= 748839539;
assign addr[11016]= 676689746;
assign addr[11017]= 603681519;
assign addr[11018]= 529907477;
assign addr[11019]= 455461206;
assign addr[11020]= 380437148;
assign addr[11021]= 304930476;
assign addr[11022]= 229036977;
assign addr[11023]= 152852926;
assign addr[11024]= 76474970;
assign addr[11025]= 0;
assign addr[11026]= -76474970;
assign addr[11027]= -152852926;
assign addr[11028]= -229036977;
assign addr[11029]= -304930476;
assign addr[11030]= -380437148;
assign addr[11031]= -455461206;
assign addr[11032]= -529907477;
assign addr[11033]= -603681519;
assign addr[11034]= -676689746;
assign addr[11035]= -748839539;
assign addr[11036]= -820039373;
assign addr[11037]= -890198924;
assign addr[11038]= -959229189;
assign addr[11039]= -1027042599;
assign addr[11040]= -1093553126;
assign addr[11041]= -1158676398;
assign addr[11042]= -1222329801;
assign addr[11043]= -1284432584;
assign addr[11044]= -1344905966;
assign addr[11045]= -1403673233;
assign addr[11046]= -1460659832;
assign addr[11047]= -1515793473;
assign addr[11048]= -1569004214;
assign addr[11049]= -1620224553;
assign addr[11050]= -1669389513;
assign addr[11051]= -1716436725;
assign addr[11052]= -1761306505;
assign addr[11053]= -1803941934;
assign addr[11054]= -1844288924;
assign addr[11055]= -1882296293;
assign addr[11056]= -1917915825;
assign addr[11057]= -1951102334;
assign addr[11058]= -1981813720;
assign addr[11059]= -2010011024;
assign addr[11060]= -2035658475;
assign addr[11061]= -2058723538;
assign addr[11062]= -2079176953;
assign addr[11063]= -2096992772;
assign addr[11064]= -2112148396;
assign addr[11065]= -2124624598;
assign addr[11066]= -2134405552;
assign addr[11067]= -2141478848;
assign addr[11068]= -2145835515;
assign addr[11069]= -2147470025;
assign addr[11070]= -2146380306;
assign addr[11071]= -2142567738;
assign addr[11072]= -2136037160;
assign addr[11073]= -2126796855;
assign addr[11074]= -2114858546;
assign addr[11075]= -2100237377;
assign addr[11076]= -2082951896;
assign addr[11077]= -2063024031;
assign addr[11078]= -2040479063;
assign addr[11079]= -2015345591;
assign addr[11080]= -1987655498;
assign addr[11081]= -1957443913;
assign addr[11082]= -1924749160;
assign addr[11083]= -1889612716;
assign addr[11084]= -1852079154;
assign addr[11085]= -1812196087;
assign addr[11086]= -1770014111;
assign addr[11087]= -1725586737;
assign addr[11088]= -1678970324;
assign addr[11089]= -1630224009;
assign addr[11090]= -1579409630;
assign addr[11091]= -1526591649;
assign addr[11092]= -1471837070;
assign addr[11093]= -1415215352;
assign addr[11094]= -1356798326;
assign addr[11095]= -1296660098;
assign addr[11096]= -1234876957;
assign addr[11097]= -1171527280;
assign addr[11098]= -1106691431;
assign addr[11099]= -1040451659;
assign addr[11100]= -972891995;
assign addr[11101]= -904098143;
assign addr[11102]= -834157373;
assign addr[11103]= -763158411;
assign addr[11104]= -691191324;
assign addr[11105]= -618347408;
assign addr[11106]= -544719071;
assign addr[11107]= -470399716;
assign addr[11108]= -395483624;
assign addr[11109]= -320065829;
assign addr[11110]= -244242007;
assign addr[11111]= -168108346;
assign addr[11112]= -91761426;
assign addr[11113]= -15298099;
assign addr[11114]= 61184634;
assign addr[11115]= 137589750;
assign addr[11116]= 213820322;
assign addr[11117]= 289779648;
assign addr[11118]= 365371365;
assign addr[11119]= 440499581;
assign addr[11120]= 515068990;
assign addr[11121]= 588984994;
assign addr[11122]= 662153826;
assign addr[11123]= 734482665;
assign addr[11124]= 805879757;
assign addr[11125]= 876254528;
assign addr[11126]= 945517704;
assign addr[11127]= 1013581418;
assign addr[11128]= 1080359326;
assign addr[11129]= 1145766716;
assign addr[11130]= 1209720613;
assign addr[11131]= 1272139887;
assign addr[11132]= 1332945355;
assign addr[11133]= 1392059879;
assign addr[11134]= 1449408469;
assign addr[11135]= 1504918373;
assign addr[11136]= 1558519173;
assign addr[11137]= 1610142873;
assign addr[11138]= 1659723983;
assign addr[11139]= 1707199606;
assign addr[11140]= 1752509516;
assign addr[11141]= 1795596234;
assign addr[11142]= 1836405100;
assign addr[11143]= 1874884346;
assign addr[11144]= 1910985158;
assign addr[11145]= 1944661739;
assign addr[11146]= 1975871368;
assign addr[11147]= 2004574453;
assign addr[11148]= 2030734582;
assign addr[11149]= 2054318569;
assign addr[11150]= 2075296495;
assign addr[11151]= 2093641749;
assign addr[11152]= 2109331059;
assign addr[11153]= 2122344521;
assign addr[11154]= 2132665626;
assign addr[11155]= 2140281282;
assign addr[11156]= 2145181827;
assign addr[11157]= 2147361045;
assign addr[11158]= 2146816171;
assign addr[11159]= 2143547897;
assign addr[11160]= 2137560369;
assign addr[11161]= 2128861181;
assign addr[11162]= 2117461370;
assign addr[11163]= 2103375398;
assign addr[11164]= 2086621133;
assign addr[11165]= 2067219829;
assign addr[11166]= 2045196100;
assign addr[11167]= 2020577882;
assign addr[11168]= 1993396407;
assign addr[11169]= 1963686155;
assign addr[11170]= 1931484818;
assign addr[11171]= 1896833245;
assign addr[11172]= 1859775393;
assign addr[11173]= 1820358275;
assign addr[11174]= 1778631892;
assign addr[11175]= 1734649179;
assign addr[11176]= 1688465931;
assign addr[11177]= 1640140734;
assign addr[11178]= 1589734894;
assign addr[11179]= 1537312353;
assign addr[11180]= 1482939614;
assign addr[11181]= 1426685652;
assign addr[11182]= 1368621831;
assign addr[11183]= 1308821808;
assign addr[11184]= 1247361445;
assign addr[11185]= 1184318708;
assign addr[11186]= 1119773573;
assign addr[11187]= 1053807919;
assign addr[11188]= 986505429;
assign addr[11189]= 917951481;
assign addr[11190]= 848233042;
assign addr[11191]= 777438554;
assign addr[11192]= 705657826;
assign addr[11193]= 632981917;
assign addr[11194]= 559503022;
assign addr[11195]= 485314355;
assign addr[11196]= 410510029;
assign addr[11197]= 335184940;
assign addr[11198]= 259434643;
assign addr[11199]= 183355234;
assign addr[11200]= 107043224;
assign addr[11201]= 30595422;
assign addr[11202]= -45891193;
assign addr[11203]= -122319591;
assign addr[11204]= -198592817;
assign addr[11205]= -274614114;
assign addr[11206]= -350287041;
assign addr[11207]= -425515602;
assign addr[11208]= -500204365;
assign addr[11209]= -574258580;
assign addr[11210]= -647584304;
assign addr[11211]= -720088517;
assign addr[11212]= -791679244;
assign addr[11213]= -862265664;
assign addr[11214]= -931758235;
assign addr[11215]= -1000068799;
assign addr[11216]= -1067110699;
assign addr[11217]= -1132798888;
assign addr[11218]= -1197050035;
assign addr[11219]= -1259782632;
assign addr[11220]= -1320917099;
assign addr[11221]= -1380375881;
assign addr[11222]= -1438083551;
assign addr[11223]= -1493966902;
assign addr[11224]= -1547955041;
assign addr[11225]= -1599979481;
assign addr[11226]= -1649974225;
assign addr[11227]= -1697875851;
assign addr[11228]= -1743623590;
assign addr[11229]= -1787159411;
assign addr[11230]= -1828428082;
assign addr[11231]= -1867377253;
assign addr[11232]= -1903957513;
assign addr[11233]= -1938122457;
assign addr[11234]= -1969828744;
assign addr[11235]= -1999036154;
assign addr[11236]= -2025707632;
assign addr[11237]= -2049809346;
assign addr[11238]= -2071310720;
assign addr[11239]= -2090184478;
assign addr[11240]= -2106406677;
assign addr[11241]= -2119956737;
assign addr[11242]= -2130817471;
assign addr[11243]= -2138975100;
assign addr[11244]= -2144419275;
assign addr[11245]= -2147143090;
assign addr[11246]= -2147143090;
assign addr[11247]= -2144419275;
assign addr[11248]= -2138975100;
assign addr[11249]= -2130817471;
assign addr[11250]= -2119956737;
assign addr[11251]= -2106406677;
assign addr[11252]= -2090184478;
assign addr[11253]= -2071310720;
assign addr[11254]= -2049809346;
assign addr[11255]= -2025707632;
assign addr[11256]= -1999036154;
assign addr[11257]= -1969828744;
assign addr[11258]= -1938122457;
assign addr[11259]= -1903957513;
assign addr[11260]= -1867377253;
assign addr[11261]= -1828428082;
assign addr[11262]= -1787159411;
assign addr[11263]= -1743623590;
assign addr[11264]= -1697875851;
assign addr[11265]= -1649974225;
assign addr[11266]= -1599979481;
assign addr[11267]= -1547955041;
assign addr[11268]= -1493966902;
assign addr[11269]= -1438083551;
assign addr[11270]= -1380375881;
assign addr[11271]= -1320917099;
assign addr[11272]= -1259782632;
assign addr[11273]= -1197050035;
assign addr[11274]= -1132798888;
assign addr[11275]= -1067110699;
assign addr[11276]= -1000068799;
assign addr[11277]= -931758235;
assign addr[11278]= -862265664;
assign addr[11279]= -791679244;
assign addr[11280]= -720088517;
assign addr[11281]= -647584304;
assign addr[11282]= -574258580;
assign addr[11283]= -500204365;
assign addr[11284]= -425515602;
assign addr[11285]= -350287041;
assign addr[11286]= -274614114;
assign addr[11287]= -198592817;
assign addr[11288]= -122319591;
assign addr[11289]= -45891193;
assign addr[11290]= 30595422;
assign addr[11291]= 107043224;
assign addr[11292]= 183355234;
assign addr[11293]= 259434643;
assign addr[11294]= 335184940;
assign addr[11295]= 410510029;
assign addr[11296]= 485314355;
assign addr[11297]= 559503022;
assign addr[11298]= 632981917;
assign addr[11299]= 705657826;
assign addr[11300]= 777438554;
assign addr[11301]= 848233042;
assign addr[11302]= 917951481;
assign addr[11303]= 986505429;
assign addr[11304]= 1053807919;
assign addr[11305]= 1119773573;
assign addr[11306]= 1184318708;
assign addr[11307]= 1247361445;
assign addr[11308]= 1308821808;
assign addr[11309]= 1368621831;
assign addr[11310]= 1426685652;
assign addr[11311]= 1482939614;
assign addr[11312]= 1537312353;
assign addr[11313]= 1589734894;
assign addr[11314]= 1640140734;
assign addr[11315]= 1688465931;
assign addr[11316]= 1734649179;
assign addr[11317]= 1778631892;
assign addr[11318]= 1820358275;
assign addr[11319]= 1859775393;
assign addr[11320]= 1896833245;
assign addr[11321]= 1931484818;
assign addr[11322]= 1963686155;
assign addr[11323]= 1993396407;
assign addr[11324]= 2020577882;
assign addr[11325]= 2045196100;
assign addr[11326]= 2067219829;
assign addr[11327]= 2086621133;
assign addr[11328]= 2103375398;
assign addr[11329]= 2117461370;
assign addr[11330]= 2128861181;
assign addr[11331]= 2137560369;
assign addr[11332]= 2143547897;
assign addr[11333]= 2146816171;
assign addr[11334]= 2147361045;
assign addr[11335]= 2145181827;
assign addr[11336]= 2140281282;
assign addr[11337]= 2132665626;
assign addr[11338]= 2122344521;
assign addr[11339]= 2109331059;
assign addr[11340]= 2093641749;
assign addr[11341]= 2075296495;
assign addr[11342]= 2054318569;
assign addr[11343]= 2030734582;
assign addr[11344]= 2004574453;
assign addr[11345]= 1975871368;
assign addr[11346]= 1944661739;
assign addr[11347]= 1910985158;
assign addr[11348]= 1874884346;
assign addr[11349]= 1836405100;
assign addr[11350]= 1795596234;
assign addr[11351]= 1752509516;
assign addr[11352]= 1707199606;
assign addr[11353]= 1659723983;
assign addr[11354]= 1610142873;
assign addr[11355]= 1558519173;
assign addr[11356]= 1504918373;
assign addr[11357]= 1449408469;
assign addr[11358]= 1392059879;
assign addr[11359]= 1332945355;
assign addr[11360]= 1272139887;
assign addr[11361]= 1209720613;
assign addr[11362]= 1145766716;
assign addr[11363]= 1080359326;
assign addr[11364]= 1013581418;
assign addr[11365]= 945517704;
assign addr[11366]= 876254528;
assign addr[11367]= 805879757;
assign addr[11368]= 734482665;
assign addr[11369]= 662153826;
assign addr[11370]= 588984994;
assign addr[11371]= 515068990;
assign addr[11372]= 440499581;
assign addr[11373]= 365371365;
assign addr[11374]= 289779648;
assign addr[11375]= 213820322;
assign addr[11376]= 137589750;
assign addr[11377]= 61184634;
assign addr[11378]= -15298099;
assign addr[11379]= -91761426;
assign addr[11380]= -168108346;
assign addr[11381]= -244242007;
assign addr[11382]= -320065829;
assign addr[11383]= -395483624;
assign addr[11384]= -470399716;
assign addr[11385]= -544719071;
assign addr[11386]= -618347408;
assign addr[11387]= -691191324;
assign addr[11388]= -763158411;
assign addr[11389]= -834157373;
assign addr[11390]= -904098143;
assign addr[11391]= -972891995;
assign addr[11392]= -1040451659;
assign addr[11393]= -1106691431;
assign addr[11394]= -1171527280;
assign addr[11395]= -1234876957;
assign addr[11396]= -1296660098;
assign addr[11397]= -1356798326;
assign addr[11398]= -1415215352;
assign addr[11399]= -1471837070;
assign addr[11400]= -1526591649;
assign addr[11401]= -1579409630;
assign addr[11402]= -1630224009;
assign addr[11403]= -1678970324;
assign addr[11404]= -1725586737;
assign addr[11405]= -1770014111;
assign addr[11406]= -1812196087;
assign addr[11407]= -1852079154;
assign addr[11408]= -1889612716;
assign addr[11409]= -1924749160;
assign addr[11410]= -1957443913;
assign addr[11411]= -1987655498;
assign addr[11412]= -2015345591;
assign addr[11413]= -2040479063;
assign addr[11414]= -2063024031;
assign addr[11415]= -2082951896;
assign addr[11416]= -2100237377;
assign addr[11417]= -2114858546;
assign addr[11418]= -2126796855;
assign addr[11419]= -2136037160;
assign addr[11420]= -2142567738;
assign addr[11421]= -2146380306;
assign addr[11422]= -2147470025;
assign addr[11423]= -2145835515;
assign addr[11424]= -2141478848;
assign addr[11425]= -2134405552;
assign addr[11426]= -2124624598;
assign addr[11427]= -2112148396;
assign addr[11428]= -2096992772;
assign addr[11429]= -2079176953;
assign addr[11430]= -2058723538;
assign addr[11431]= -2035658475;
assign addr[11432]= -2010011024;
assign addr[11433]= -1981813720;
assign addr[11434]= -1951102334;
assign addr[11435]= -1917915825;
assign addr[11436]= -1882296293;
assign addr[11437]= -1844288924;
assign addr[11438]= -1803941934;
assign addr[11439]= -1761306505;
assign addr[11440]= -1716436725;
assign addr[11441]= -1669389513;
assign addr[11442]= -1620224553;
assign addr[11443]= -1569004214;
assign addr[11444]= -1515793473;
assign addr[11445]= -1460659832;
assign addr[11446]= -1403673233;
assign addr[11447]= -1344905966;
assign addr[11448]= -1284432584;
assign addr[11449]= -1222329801;
assign addr[11450]= -1158676398;
assign addr[11451]= -1093553126;
assign addr[11452]= -1027042599;
assign addr[11453]= -959229189;
assign addr[11454]= -890198924;
assign addr[11455]= -820039373;
assign addr[11456]= -748839539;
assign addr[11457]= -676689746;
assign addr[11458]= -603681519;
assign addr[11459]= -529907477;
assign addr[11460]= -455461206;
assign addr[11461]= -380437148;
assign addr[11462]= -304930476;
assign addr[11463]= -229036977;
assign addr[11464]= -152852926;
assign addr[11465]= -76474970;
assign addr[11466]= 0;
assign addr[11467]= 76474970;
assign addr[11468]= 152852926;
assign addr[11469]= 229036977;
assign addr[11470]= 304930476;
assign addr[11471]= 380437148;
assign addr[11472]= 455461206;
assign addr[11473]= 529907477;
assign addr[11474]= 603681519;
assign addr[11475]= 676689746;
assign addr[11476]= 748839539;
assign addr[11477]= 820039373;
assign addr[11478]= 890198924;
assign addr[11479]= 959229189;
assign addr[11480]= 1027042599;
assign addr[11481]= 1093553126;
assign addr[11482]= 1158676398;
assign addr[11483]= 1222329801;
assign addr[11484]= 1284432584;
assign addr[11485]= 1344905966;
assign addr[11486]= 1403673233;
assign addr[11487]= 1460659832;
assign addr[11488]= 1515793473;
assign addr[11489]= 1569004214;
assign addr[11490]= 1620224553;
assign addr[11491]= 1669389513;
assign addr[11492]= 1716436725;
assign addr[11493]= 1761306505;
assign addr[11494]= 1803941934;
assign addr[11495]= 1844288924;
assign addr[11496]= 1882296293;
assign addr[11497]= 1917915825;
assign addr[11498]= 1951102334;
assign addr[11499]= 1981813720;
assign addr[11500]= 2010011024;
assign addr[11501]= 2035658475;
assign addr[11502]= 2058723538;
assign addr[11503]= 2079176953;
assign addr[11504]= 2096992772;
assign addr[11505]= 2112148396;
assign addr[11506]= 2124624598;
assign addr[11507]= 2134405552;
assign addr[11508]= 2141478848;
assign addr[11509]= 2145835515;
assign addr[11510]= 2147470025;
assign addr[11511]= 2146380306;
assign addr[11512]= 2142567738;
assign addr[11513]= 2136037160;
assign addr[11514]= 2126796855;
assign addr[11515]= 2114858546;
assign addr[11516]= 2100237377;
assign addr[11517]= 2082951896;
assign addr[11518]= 2063024031;
assign addr[11519]= 2040479063;
assign addr[11520]= 2015345591;
assign addr[11521]= 1987655498;
assign addr[11522]= 1957443913;
assign addr[11523]= 1924749160;
assign addr[11524]= 1889612716;
assign addr[11525]= 1852079154;
assign addr[11526]= 1812196087;
assign addr[11527]= 1770014111;
assign addr[11528]= 1725586737;
assign addr[11529]= 1678970324;
assign addr[11530]= 1630224009;
assign addr[11531]= 1579409630;
assign addr[11532]= 1526591649;
assign addr[11533]= 1471837070;
assign addr[11534]= 1415215352;
assign addr[11535]= 1356798326;
assign addr[11536]= 1296660098;
assign addr[11537]= 1234876957;
assign addr[11538]= 1171527280;
assign addr[11539]= 1106691431;
assign addr[11540]= 1040451659;
assign addr[11541]= 972891995;
assign addr[11542]= 904098143;
assign addr[11543]= 834157373;
assign addr[11544]= 763158411;
assign addr[11545]= 691191324;
assign addr[11546]= 618347408;
assign addr[11547]= 544719071;
assign addr[11548]= 470399716;
assign addr[11549]= 395483624;
assign addr[11550]= 320065829;
assign addr[11551]= 244242007;
assign addr[11552]= 168108346;
assign addr[11553]= 91761426;
assign addr[11554]= 15298099;
assign addr[11555]= -61184634;
assign addr[11556]= -137589750;
assign addr[11557]= -213820322;
assign addr[11558]= -289779648;
assign addr[11559]= -365371365;
assign addr[11560]= -440499581;
assign addr[11561]= -515068990;
assign addr[11562]= -588984994;
assign addr[11563]= -662153826;
assign addr[11564]= -734482665;
assign addr[11565]= -805879757;
assign addr[11566]= -876254528;
assign addr[11567]= -945517704;
assign addr[11568]= -1013581418;
assign addr[11569]= -1080359326;
assign addr[11570]= -1145766716;
assign addr[11571]= -1209720613;
assign addr[11572]= -1272139887;
assign addr[11573]= -1332945355;
assign addr[11574]= -1392059879;
assign addr[11575]= -1449408469;
assign addr[11576]= -1504918373;
assign addr[11577]= -1558519173;
assign addr[11578]= -1610142873;
assign addr[11579]= -1659723983;
assign addr[11580]= -1707199606;
assign addr[11581]= -1752509516;
assign addr[11582]= -1795596234;
assign addr[11583]= -1836405100;
assign addr[11584]= -1874884346;
assign addr[11585]= -1910985158;
assign addr[11586]= -1944661739;
assign addr[11587]= -1975871368;
assign addr[11588]= -2004574453;
assign addr[11589]= -2030734582;
assign addr[11590]= -2054318569;
assign addr[11591]= -2075296495;
assign addr[11592]= -2093641749;
assign addr[11593]= -2109331059;
assign addr[11594]= -2122344521;
assign addr[11595]= -2132665626;
assign addr[11596]= -2140281282;
assign addr[11597]= -2145181827;
assign addr[11598]= -2147361045;
assign addr[11599]= -2146816171;
assign addr[11600]= -2143547897;
assign addr[11601]= -2137560369;
assign addr[11602]= -2128861181;
assign addr[11603]= -2117461370;
assign addr[11604]= -2103375398;
assign addr[11605]= -2086621133;
assign addr[11606]= -2067219829;
assign addr[11607]= -2045196100;
assign addr[11608]= -2020577882;
assign addr[11609]= -1993396407;
assign addr[11610]= -1963686155;
assign addr[11611]= -1931484818;
assign addr[11612]= -1896833245;
assign addr[11613]= -1859775393;
assign addr[11614]= -1820358275;
assign addr[11615]= -1778631892;
assign addr[11616]= -1734649179;
assign addr[11617]= -1688465931;
assign addr[11618]= -1640140734;
assign addr[11619]= -1589734894;
assign addr[11620]= -1537312353;
assign addr[11621]= -1482939614;
assign addr[11622]= -1426685652;
assign addr[11623]= -1368621831;
assign addr[11624]= -1308821808;
assign addr[11625]= -1247361445;
assign addr[11626]= -1184318708;
assign addr[11627]= -1119773573;
assign addr[11628]= -1053807919;
assign addr[11629]= -986505429;
assign addr[11630]= -917951481;
assign addr[11631]= -848233042;
assign addr[11632]= -777438554;
assign addr[11633]= -705657826;
assign addr[11634]= -632981917;
assign addr[11635]= -559503022;
assign addr[11636]= -485314355;
assign addr[11637]= -410510029;
assign addr[11638]= -335184940;
assign addr[11639]= -259434643;
assign addr[11640]= -183355234;
assign addr[11641]= -107043224;
assign addr[11642]= -30595422;
assign addr[11643]= 45891193;
assign addr[11644]= 122319591;
assign addr[11645]= 198592817;
assign addr[11646]= 274614114;
assign addr[11647]= 350287041;
assign addr[11648]= 425515602;
assign addr[11649]= 500204365;
assign addr[11650]= 574258580;
assign addr[11651]= 647584304;
assign addr[11652]= 720088517;
assign addr[11653]= 791679244;
assign addr[11654]= 862265664;
assign addr[11655]= 931758235;
assign addr[11656]= 1000068799;
assign addr[11657]= 1067110699;
assign addr[11658]= 1132798888;
assign addr[11659]= 1197050035;
assign addr[11660]= 1259782632;
assign addr[11661]= 1320917099;
assign addr[11662]= 1380375881;
assign addr[11663]= 1438083551;
assign addr[11664]= 1493966902;
assign addr[11665]= 1547955041;
assign addr[11666]= 1599979481;
assign addr[11667]= 1649974225;
assign addr[11668]= 1697875851;
assign addr[11669]= 1743623590;
assign addr[11670]= 1787159411;
assign addr[11671]= 1828428082;
assign addr[11672]= 1867377253;
assign addr[11673]= 1903957513;
assign addr[11674]= 1938122457;
assign addr[11675]= 1969828744;
assign addr[11676]= 1999036154;
assign addr[11677]= 2025707632;
assign addr[11678]= 2049809346;
assign addr[11679]= 2071310720;
assign addr[11680]= 2090184478;
assign addr[11681]= 2106406677;
assign addr[11682]= 2119956737;
assign addr[11683]= 2130817471;
assign addr[11684]= 2138975100;
assign addr[11685]= 2144419275;
assign addr[11686]= 2147143090;
assign addr[11687]= 2147143090;
assign addr[11688]= 2144419275;
assign addr[11689]= 2138975100;
assign addr[11690]= 2130817471;
assign addr[11691]= 2119956737;
assign addr[11692]= 2106406677;
assign addr[11693]= 2090184478;
assign addr[11694]= 2071310720;
assign addr[11695]= 2049809346;
assign addr[11696]= 2025707632;
assign addr[11697]= 1999036154;
assign addr[11698]= 1969828744;
assign addr[11699]= 1938122457;
assign addr[11700]= 1903957513;
assign addr[11701]= 1867377253;
assign addr[11702]= 1828428082;
assign addr[11703]= 1787159411;
assign addr[11704]= 1743623590;
assign addr[11705]= 1697875851;
assign addr[11706]= 1649974225;
assign addr[11707]= 1599979481;
assign addr[11708]= 1547955041;
assign addr[11709]= 1493966902;
assign addr[11710]= 1438083551;
assign addr[11711]= 1380375881;
assign addr[11712]= 1320917099;
assign addr[11713]= 1259782632;
assign addr[11714]= 1197050035;
assign addr[11715]= 1132798888;
assign addr[11716]= 1067110699;
assign addr[11717]= 1000068799;
assign addr[11718]= 931758235;
assign addr[11719]= 862265664;
assign addr[11720]= 791679244;
assign addr[11721]= 720088517;
assign addr[11722]= 647584304;
assign addr[11723]= 574258580;
assign addr[11724]= 500204365;
assign addr[11725]= 425515602;
assign addr[11726]= 350287041;
assign addr[11727]= 274614114;
assign addr[11728]= 198592817;
assign addr[11729]= 122319591;
assign addr[11730]= 45891193;
assign addr[11731]= -30595422;
assign addr[11732]= -107043224;
assign addr[11733]= -183355234;
assign addr[11734]= -259434643;
assign addr[11735]= -335184940;
assign addr[11736]= -410510029;
assign addr[11737]= -485314355;
assign addr[11738]= -559503022;
assign addr[11739]= -632981917;
assign addr[11740]= -705657826;
assign addr[11741]= -777438554;
assign addr[11742]= -848233042;
assign addr[11743]= -917951481;
assign addr[11744]= -986505429;
assign addr[11745]= -1053807919;
assign addr[11746]= -1119773573;
assign addr[11747]= -1184318708;
assign addr[11748]= -1247361445;
assign addr[11749]= -1308821808;
assign addr[11750]= -1368621831;
assign addr[11751]= -1426685652;
assign addr[11752]= -1482939614;
assign addr[11753]= -1537312353;
assign addr[11754]= -1589734894;
assign addr[11755]= -1640140734;
assign addr[11756]= -1688465931;
assign addr[11757]= -1734649179;
assign addr[11758]= -1778631892;
assign addr[11759]= -1820358275;
assign addr[11760]= -1859775393;
assign addr[11761]= -1896833245;
assign addr[11762]= -1931484818;
assign addr[11763]= -1963686155;
assign addr[11764]= -1993396407;
assign addr[11765]= -2020577882;
assign addr[11766]= -2045196100;
assign addr[11767]= -2067219829;
assign addr[11768]= -2086621133;
assign addr[11769]= -2103375398;
assign addr[11770]= -2117461370;
assign addr[11771]= -2128861181;
assign addr[11772]= -2137560369;
assign addr[11773]= -2143547897;
assign addr[11774]= -2146816171;
assign addr[11775]= -2147361045;
assign addr[11776]= -2145181827;
assign addr[11777]= -2140281282;
assign addr[11778]= -2132665626;
assign addr[11779]= -2122344521;
assign addr[11780]= -2109331059;
assign addr[11781]= -2093641749;
assign addr[11782]= -2075296495;
assign addr[11783]= -2054318569;
assign addr[11784]= -2030734582;
assign addr[11785]= -2004574453;
assign addr[11786]= -1975871368;
assign addr[11787]= -1944661739;
assign addr[11788]= -1910985158;
assign addr[11789]= -1874884346;
assign addr[11790]= -1836405100;
assign addr[11791]= -1795596234;
assign addr[11792]= -1752509516;
assign addr[11793]= -1707199606;
assign addr[11794]= -1659723983;
assign addr[11795]= -1610142873;
assign addr[11796]= -1558519173;
assign addr[11797]= -1504918373;
assign addr[11798]= -1449408469;
assign addr[11799]= -1392059879;
assign addr[11800]= -1332945355;
assign addr[11801]= -1272139887;
assign addr[11802]= -1209720613;
assign addr[11803]= -1145766716;
assign addr[11804]= -1080359326;
assign addr[11805]= -1013581418;
assign addr[11806]= -945517704;
assign addr[11807]= -876254528;
assign addr[11808]= -805879757;
assign addr[11809]= -734482665;
assign addr[11810]= -662153826;
assign addr[11811]= -588984994;
assign addr[11812]= -515068990;
assign addr[11813]= -440499581;
assign addr[11814]= -365371365;
assign addr[11815]= -289779648;
assign addr[11816]= -213820322;
assign addr[11817]= -137589750;
assign addr[11818]= -61184634;
assign addr[11819]= 15298099;
assign addr[11820]= 91761426;
assign addr[11821]= 168108346;
assign addr[11822]= 244242007;
assign addr[11823]= 320065829;
assign addr[11824]= 395483624;
assign addr[11825]= 470399716;
assign addr[11826]= 544719071;
assign addr[11827]= 618347408;
assign addr[11828]= 691191324;
assign addr[11829]= 763158411;
assign addr[11830]= 834157373;
assign addr[11831]= 904098143;
assign addr[11832]= 972891995;
assign addr[11833]= 1040451659;
assign addr[11834]= 1106691431;
assign addr[11835]= 1171527280;
assign addr[11836]= 1234876957;
assign addr[11837]= 1296660098;
assign addr[11838]= 1356798326;
assign addr[11839]= 1415215352;
assign addr[11840]= 1471837070;
assign addr[11841]= 1526591649;
assign addr[11842]= 1579409630;
assign addr[11843]= 1630224009;
assign addr[11844]= 1678970324;
assign addr[11845]= 1725586737;
assign addr[11846]= 1770014111;
assign addr[11847]= 1812196087;
assign addr[11848]= 1852079154;
assign addr[11849]= 1889612716;
assign addr[11850]= 1924749160;
assign addr[11851]= 1957443913;
assign addr[11852]= 1987655498;
assign addr[11853]= 2015345591;
assign addr[11854]= 2040479063;
assign addr[11855]= 2063024031;
assign addr[11856]= 2082951896;
assign addr[11857]= 2100237377;
assign addr[11858]= 2114858546;
assign addr[11859]= 2126796855;
assign addr[11860]= 2136037160;
assign addr[11861]= 2142567738;
assign addr[11862]= 2146380306;
assign addr[11863]= 2147470025;
assign addr[11864]= 2145835515;
assign addr[11865]= 2141478848;
assign addr[11866]= 2134405552;
assign addr[11867]= 2124624598;
assign addr[11868]= 2112148396;
assign addr[11869]= 2096992772;
assign addr[11870]= 2079176953;
assign addr[11871]= 2058723538;
assign addr[11872]= 2035658475;
assign addr[11873]= 2010011024;
assign addr[11874]= 1981813720;
assign addr[11875]= 1951102334;
assign addr[11876]= 1917915825;
assign addr[11877]= 1882296293;
assign addr[11878]= 1844288924;
assign addr[11879]= 1803941934;
assign addr[11880]= 1761306505;
assign addr[11881]= 1716436725;
assign addr[11882]= 1669389513;
assign addr[11883]= 1620224553;
assign addr[11884]= 1569004214;
assign addr[11885]= 1515793473;
assign addr[11886]= 1460659832;
assign addr[11887]= 1403673233;
assign addr[11888]= 1344905966;
assign addr[11889]= 1284432584;
assign addr[11890]= 1222329801;
assign addr[11891]= 1158676398;
assign addr[11892]= 1093553126;
assign addr[11893]= 1027042599;
assign addr[11894]= 959229189;
assign addr[11895]= 890198924;
assign addr[11896]= 820039373;
assign addr[11897]= 748839539;
assign addr[11898]= 676689746;
assign addr[11899]= 603681519;
assign addr[11900]= 529907477;
assign addr[11901]= 455461206;
assign addr[11902]= 380437148;
assign addr[11903]= 304930476;
assign addr[11904]= 229036977;
assign addr[11905]= 152852926;
assign addr[11906]= 76474970;
assign addr[11907]= 0;
assign addr[11908]= -76474970;
assign addr[11909]= -152852926;
assign addr[11910]= -229036977;
assign addr[11911]= -304930476;
assign addr[11912]= -380437148;
assign addr[11913]= -455461206;
assign addr[11914]= -529907477;
assign addr[11915]= -603681519;
assign addr[11916]= -676689746;
assign addr[11917]= -748839539;
assign addr[11918]= -820039373;
assign addr[11919]= -890198924;
assign addr[11920]= -959229189;
assign addr[11921]= -1027042599;
assign addr[11922]= -1093553126;
assign addr[11923]= -1158676398;
assign addr[11924]= -1222329801;
assign addr[11925]= -1284432584;
assign addr[11926]= -1344905966;
assign addr[11927]= -1403673233;
assign addr[11928]= -1460659832;
assign addr[11929]= -1515793473;
assign addr[11930]= -1569004214;
assign addr[11931]= -1620224553;
assign addr[11932]= -1669389513;
assign addr[11933]= -1716436725;
assign addr[11934]= -1761306505;
assign addr[11935]= -1803941934;
assign addr[11936]= -1844288924;
assign addr[11937]= -1882296293;
assign addr[11938]= -1917915825;
assign addr[11939]= -1951102334;
assign addr[11940]= -1981813720;
assign addr[11941]= -2010011024;
assign addr[11942]= -2035658475;
assign addr[11943]= -2058723538;
assign addr[11944]= -2079176953;
assign addr[11945]= -2096992772;
assign addr[11946]= -2112148396;
assign addr[11947]= -2124624598;
assign addr[11948]= -2134405552;
assign addr[11949]= -2141478848;
assign addr[11950]= -2145835515;
assign addr[11951]= -2147470025;
assign addr[11952]= -2146380306;
assign addr[11953]= -2142567738;
assign addr[11954]= -2136037160;
assign addr[11955]= -2126796855;
assign addr[11956]= -2114858546;
assign addr[11957]= -2100237377;
assign addr[11958]= -2082951896;
assign addr[11959]= -2063024031;
assign addr[11960]= -2040479063;
assign addr[11961]= -2015345591;
assign addr[11962]= -1987655498;
assign addr[11963]= -1957443913;
assign addr[11964]= -1924749160;
assign addr[11965]= -1889612716;
assign addr[11966]= -1852079154;
assign addr[11967]= -1812196087;
assign addr[11968]= -1770014111;
assign addr[11969]= -1725586737;
assign addr[11970]= -1678970324;
assign addr[11971]= -1630224009;
assign addr[11972]= -1579409630;
assign addr[11973]= -1526591649;
assign addr[11974]= -1471837070;
assign addr[11975]= -1415215352;
assign addr[11976]= -1356798326;
assign addr[11977]= -1296660098;
assign addr[11978]= -1234876957;
assign addr[11979]= -1171527280;
assign addr[11980]= -1106691431;
assign addr[11981]= -1040451659;
assign addr[11982]= -972891995;
assign addr[11983]= -904098143;
assign addr[11984]= -834157373;
assign addr[11985]= -763158411;
assign addr[11986]= -691191324;
assign addr[11987]= -618347408;
assign addr[11988]= -544719071;
assign addr[11989]= -470399716;
assign addr[11990]= -395483624;
assign addr[11991]= -320065829;
assign addr[11992]= -244242007;
assign addr[11993]= -168108346;
assign addr[11994]= -91761426;
assign addr[11995]= -15298099;
assign addr[11996]= 61184634;
assign addr[11997]= 137589750;
assign addr[11998]= 213820322;
assign addr[11999]= 289779648;
assign addr[12000]= 365371365;
assign addr[12001]= 440499581;
assign addr[12002]= 515068990;
assign addr[12003]= 588984994;
assign addr[12004]= 662153826;
assign addr[12005]= 734482665;
assign addr[12006]= 805879757;
assign addr[12007]= 876254528;
assign addr[12008]= 945517704;
assign addr[12009]= 1013581418;
assign addr[12010]= 1080359326;
assign addr[12011]= 1145766716;
assign addr[12012]= 1209720613;
assign addr[12013]= 1272139887;
assign addr[12014]= 1332945355;
assign addr[12015]= 1392059879;
assign addr[12016]= 1449408469;
assign addr[12017]= 1504918373;
assign addr[12018]= 1558519173;
assign addr[12019]= 1610142873;
assign addr[12020]= 1659723983;
assign addr[12021]= 1707199606;
assign addr[12022]= 1752509516;
assign addr[12023]= 1795596234;
assign addr[12024]= 1836405100;
assign addr[12025]= 1874884346;
assign addr[12026]= 1910985158;
assign addr[12027]= 1944661739;
assign addr[12028]= 1975871368;
assign addr[12029]= 2004574453;
assign addr[12030]= 2030734582;
assign addr[12031]= 2054318569;
assign addr[12032]= 2075296495;
assign addr[12033]= 2093641749;
assign addr[12034]= 2109331059;
assign addr[12035]= 2122344521;
assign addr[12036]= 2132665626;
assign addr[12037]= 2140281282;
assign addr[12038]= 2145181827;
assign addr[12039]= 2147361045;
assign addr[12040]= 2146816171;
assign addr[12041]= 2143547897;
assign addr[12042]= 2137560369;
assign addr[12043]= 2128861181;
assign addr[12044]= 2117461370;
assign addr[12045]= 2103375398;
assign addr[12046]= 2086621133;
assign addr[12047]= 2067219829;
assign addr[12048]= 2045196100;
assign addr[12049]= 2020577882;
assign addr[12050]= 1993396407;
assign addr[12051]= 1963686155;
assign addr[12052]= 1931484818;
assign addr[12053]= 1896833245;
assign addr[12054]= 1859775393;
assign addr[12055]= 1820358275;
assign addr[12056]= 1778631892;
assign addr[12057]= 1734649179;
assign addr[12058]= 1688465931;
assign addr[12059]= 1640140734;
assign addr[12060]= 1589734894;
assign addr[12061]= 1537312353;
assign addr[12062]= 1482939614;
assign addr[12063]= 1426685652;
assign addr[12064]= 1368621831;
assign addr[12065]= 1308821808;
assign addr[12066]= 1247361445;
assign addr[12067]= 1184318708;
assign addr[12068]= 1119773573;
assign addr[12069]= 1053807919;
assign addr[12070]= 986505429;
assign addr[12071]= 917951481;
assign addr[12072]= 848233042;
assign addr[12073]= 777438554;
assign addr[12074]= 705657826;
assign addr[12075]= 632981917;
assign addr[12076]= 559503022;
assign addr[12077]= 485314355;
assign addr[12078]= 410510029;
assign addr[12079]= 335184940;
assign addr[12080]= 259434643;
assign addr[12081]= 183355234;
assign addr[12082]= 107043224;
assign addr[12083]= 30595422;
assign addr[12084]= -45891193;
assign addr[12085]= -122319591;
assign addr[12086]= -198592817;
assign addr[12087]= -274614114;
assign addr[12088]= -350287041;
assign addr[12089]= -425515602;
assign addr[12090]= -500204365;
assign addr[12091]= -574258580;
assign addr[12092]= -647584304;
assign addr[12093]= -720088517;
assign addr[12094]= -791679244;
assign addr[12095]= -862265664;
assign addr[12096]= -931758235;
assign addr[12097]= -1000068799;
assign addr[12098]= -1067110699;
assign addr[12099]= -1132798888;
assign addr[12100]= -1197050035;
assign addr[12101]= -1259782632;
assign addr[12102]= -1320917099;
assign addr[12103]= -1380375881;
assign addr[12104]= -1438083551;
assign addr[12105]= -1493966902;
assign addr[12106]= -1547955041;
assign addr[12107]= -1599979481;
assign addr[12108]= -1649974225;
assign addr[12109]= -1697875851;
assign addr[12110]= -1743623590;
assign addr[12111]= -1787159411;
assign addr[12112]= -1828428082;
assign addr[12113]= -1867377253;
assign addr[12114]= -1903957513;
assign addr[12115]= -1938122457;
assign addr[12116]= -1969828744;
assign addr[12117]= -1999036154;
assign addr[12118]= -2025707632;
assign addr[12119]= -2049809346;
assign addr[12120]= -2071310720;
assign addr[12121]= -2090184478;
assign addr[12122]= -2106406677;
assign addr[12123]= -2119956737;
assign addr[12124]= -2130817471;
assign addr[12125]= -2138975100;
assign addr[12126]= -2144419275;
assign addr[12127]= -2147143090;
assign addr[12128]= -2147143090;
assign addr[12129]= -2144419275;
assign addr[12130]= -2138975100;
assign addr[12131]= -2130817471;
assign addr[12132]= -2119956737;
assign addr[12133]= -2106406677;
assign addr[12134]= -2090184478;
assign addr[12135]= -2071310720;
assign addr[12136]= -2049809346;
assign addr[12137]= -2025707632;
assign addr[12138]= -1999036154;
assign addr[12139]= -1969828744;
assign addr[12140]= -1938122457;
assign addr[12141]= -1903957513;
assign addr[12142]= -1867377253;
assign addr[12143]= -1828428082;
assign addr[12144]= -1787159411;
assign addr[12145]= -1743623590;
assign addr[12146]= -1697875851;
assign addr[12147]= -1649974225;
assign addr[12148]= -1599979481;
assign addr[12149]= -1547955041;
assign addr[12150]= -1493966902;
assign addr[12151]= -1438083551;
assign addr[12152]= -1380375881;
assign addr[12153]= -1320917099;
assign addr[12154]= -1259782632;
assign addr[12155]= -1197050035;
assign addr[12156]= -1132798888;
assign addr[12157]= -1067110699;
assign addr[12158]= -1000068799;
assign addr[12159]= -931758235;
assign addr[12160]= -862265664;
assign addr[12161]= -791679244;
assign addr[12162]= -720088517;
assign addr[12163]= -647584304;
assign addr[12164]= -574258580;
assign addr[12165]= -500204365;
assign addr[12166]= -425515602;
assign addr[12167]= -350287041;
assign addr[12168]= -274614114;
assign addr[12169]= -198592817;
assign addr[12170]= -122319591;
assign addr[12171]= -45891193;
assign addr[12172]= 30595422;
assign addr[12173]= 107043224;
assign addr[12174]= 183355234;
assign addr[12175]= 259434643;
assign addr[12176]= 335184940;
assign addr[12177]= 410510029;
assign addr[12178]= 485314355;
assign addr[12179]= 559503022;
assign addr[12180]= 632981917;
assign addr[12181]= 705657826;
assign addr[12182]= 777438554;
assign addr[12183]= 848233042;
assign addr[12184]= 917951481;
assign addr[12185]= 986505429;
assign addr[12186]= 1053807919;
assign addr[12187]= 1119773573;
assign addr[12188]= 1184318708;
assign addr[12189]= 1247361445;
assign addr[12190]= 1308821808;
assign addr[12191]= 1368621831;
assign addr[12192]= 1426685652;
assign addr[12193]= 1482939614;
assign addr[12194]= 1537312353;
assign addr[12195]= 1589734894;
assign addr[12196]= 1640140734;
assign addr[12197]= 1688465931;
assign addr[12198]= 1734649179;
assign addr[12199]= 1778631892;
assign addr[12200]= 1820358275;
assign addr[12201]= 1859775393;
assign addr[12202]= 1896833245;
assign addr[12203]= 1931484818;
assign addr[12204]= 1963686155;
assign addr[12205]= 1993396407;
assign addr[12206]= 2020577882;
assign addr[12207]= 2045196100;
assign addr[12208]= 2067219829;
assign addr[12209]= 2086621133;
assign addr[12210]= 2103375398;
assign addr[12211]= 2117461370;
assign addr[12212]= 2128861181;
assign addr[12213]= 2137560369;
assign addr[12214]= 2143547897;
assign addr[12215]= 2146816171;
assign addr[12216]= 2147361045;
assign addr[12217]= 2145181827;
assign addr[12218]= 2140281282;
assign addr[12219]= 2132665626;
assign addr[12220]= 2122344521;
assign addr[12221]= 2109331059;
assign addr[12222]= 2093641749;
assign addr[12223]= 2075296495;
assign addr[12224]= 2054318569;
assign addr[12225]= 2030734582;
assign addr[12226]= 2004574453;
assign addr[12227]= 1975871368;
assign addr[12228]= 1944661739;
assign addr[12229]= 1910985158;
assign addr[12230]= 1874884346;
assign addr[12231]= 1836405100;
assign addr[12232]= 1795596234;
assign addr[12233]= 1752509516;
assign addr[12234]= 1707199606;
assign addr[12235]= 1659723983;
assign addr[12236]= 1610142873;
assign addr[12237]= 1558519173;
assign addr[12238]= 1504918373;
assign addr[12239]= 1449408469;
assign addr[12240]= 1392059879;
assign addr[12241]= 1332945355;
assign addr[12242]= 1272139887;
assign addr[12243]= 1209720613;
assign addr[12244]= 1145766716;
assign addr[12245]= 1080359326;
assign addr[12246]= 1013581418;
assign addr[12247]= 945517704;
assign addr[12248]= 876254528;
assign addr[12249]= 805879757;
assign addr[12250]= 734482665;
assign addr[12251]= 662153826;
assign addr[12252]= 588984994;
assign addr[12253]= 515068990;
assign addr[12254]= 440499581;
assign addr[12255]= 365371365;
assign addr[12256]= 289779648;
assign addr[12257]= 213820322;
assign addr[12258]= 137589750;
assign addr[12259]= 61184634;
assign addr[12260]= -15298099;
assign addr[12261]= -91761426;
assign addr[12262]= -168108346;
assign addr[12263]= -244242007;
assign addr[12264]= -320065829;
assign addr[12265]= -395483624;
assign addr[12266]= -470399716;
assign addr[12267]= -544719071;
assign addr[12268]= -618347408;
assign addr[12269]= -691191324;
assign addr[12270]= -763158411;
assign addr[12271]= -834157373;
assign addr[12272]= -904098143;
assign addr[12273]= -972891995;
assign addr[12274]= -1040451659;
assign addr[12275]= -1106691431;
assign addr[12276]= -1171527280;
assign addr[12277]= -1234876957;
assign addr[12278]= -1296660098;
assign addr[12279]= -1356798326;
assign addr[12280]= -1415215352;
assign addr[12281]= -1471837070;
assign addr[12282]= -1526591649;
assign addr[12283]= -1579409630;
assign addr[12284]= -1630224009;
assign addr[12285]= -1678970324;
assign addr[12286]= -1725586737;
assign addr[12287]= -1770014111;
assign addr[12288]= -1812196087;
assign addr[12289]= -1852079154;
assign addr[12290]= -1889612716;
assign addr[12291]= -1924749160;
assign addr[12292]= -1957443913;
assign addr[12293]= -1987655498;
assign addr[12294]= -2015345591;
assign addr[12295]= -2040479063;
assign addr[12296]= -2063024031;
assign addr[12297]= -2082951896;
assign addr[12298]= -2100237377;
assign addr[12299]= -2114858546;
assign addr[12300]= -2126796855;
assign addr[12301]= -2136037160;
assign addr[12302]= -2142567738;
assign addr[12303]= -2146380306;
assign addr[12304]= -2147470025;
assign addr[12305]= -2145835515;
assign addr[12306]= -2141478848;
assign addr[12307]= -2134405552;
assign addr[12308]= -2124624598;
assign addr[12309]= -2112148396;
assign addr[12310]= -2096992772;
assign addr[12311]= -2079176953;
assign addr[12312]= -2058723538;
assign addr[12313]= -2035658475;
assign addr[12314]= -2010011024;
assign addr[12315]= -1981813720;
assign addr[12316]= -1951102334;
assign addr[12317]= -1917915825;
assign addr[12318]= -1882296293;
assign addr[12319]= -1844288924;
assign addr[12320]= -1803941934;
assign addr[12321]= -1761306505;
assign addr[12322]= -1716436725;
assign addr[12323]= -1669389513;
assign addr[12324]= -1620224553;
assign addr[12325]= -1569004214;
assign addr[12326]= -1515793473;
assign addr[12327]= -1460659832;
assign addr[12328]= -1403673233;
assign addr[12329]= -1344905966;
assign addr[12330]= -1284432584;
assign addr[12331]= -1222329801;
assign addr[12332]= -1158676398;
assign addr[12333]= -1093553126;
assign addr[12334]= -1027042599;
assign addr[12335]= -959229189;
assign addr[12336]= -890198924;
assign addr[12337]= -820039373;
assign addr[12338]= -748839539;
assign addr[12339]= -676689746;
assign addr[12340]= -603681519;
assign addr[12341]= -529907477;
assign addr[12342]= -455461206;
assign addr[12343]= -380437148;
assign addr[12344]= -304930476;
assign addr[12345]= -229036977;
assign addr[12346]= -152852926;
assign addr[12347]= -76474970;
assign addr[12348]= 0;
assign addr[12349]= 76474970;
assign addr[12350]= 152852926;
assign addr[12351]= 229036977;
assign addr[12352]= 304930476;
assign addr[12353]= 380437148;
assign addr[12354]= 455461206;
assign addr[12355]= 529907477;
assign addr[12356]= 603681519;
assign addr[12357]= 676689746;
assign addr[12358]= 748839539;
assign addr[12359]= 820039373;
assign addr[12360]= 890198924;
assign addr[12361]= 959229189;
assign addr[12362]= 1027042599;
assign addr[12363]= 1093553126;
assign addr[12364]= 1158676398;
assign addr[12365]= 1222329801;
assign addr[12366]= 1284432584;
assign addr[12367]= 1344905966;
assign addr[12368]= 1403673233;
assign addr[12369]= 1460659832;
assign addr[12370]= 1515793473;
assign addr[12371]= 1569004214;
assign addr[12372]= 1620224553;
assign addr[12373]= 1669389513;
assign addr[12374]= 1716436725;
assign addr[12375]= 1761306505;
assign addr[12376]= 1803941934;
assign addr[12377]= 1844288924;
assign addr[12378]= 1882296293;
assign addr[12379]= 1917915825;
assign addr[12380]= 1951102334;
assign addr[12381]= 1981813720;
assign addr[12382]= 2010011024;
assign addr[12383]= 2035658475;
assign addr[12384]= 2058723538;
assign addr[12385]= 2079176953;
assign addr[12386]= 2096992772;
assign addr[12387]= 2112148396;
assign addr[12388]= 2124624598;
assign addr[12389]= 2134405552;
assign addr[12390]= 2141478848;
assign addr[12391]= 2145835515;
assign addr[12392]= 2147470025;
assign addr[12393]= 2146380306;
assign addr[12394]= 2142567738;
assign addr[12395]= 2136037160;
assign addr[12396]= 2126796855;
assign addr[12397]= 2114858546;
assign addr[12398]= 2100237377;
assign addr[12399]= 2082951896;
assign addr[12400]= 2063024031;
assign addr[12401]= 2040479063;
assign addr[12402]= 2015345591;
assign addr[12403]= 1987655498;
assign addr[12404]= 1957443913;
assign addr[12405]= 1924749160;
assign addr[12406]= 1889612716;
assign addr[12407]= 1852079154;
assign addr[12408]= 1812196087;
assign addr[12409]= 1770014111;
assign addr[12410]= 1725586737;
assign addr[12411]= 1678970324;
assign addr[12412]= 1630224009;
assign addr[12413]= 1579409630;
assign addr[12414]= 1526591649;
assign addr[12415]= 1471837070;
assign addr[12416]= 1415215352;
assign addr[12417]= 1356798326;
assign addr[12418]= 1296660098;
assign addr[12419]= 1234876957;
assign addr[12420]= 1171527280;
assign addr[12421]= 1106691431;
assign addr[12422]= 1040451659;
assign addr[12423]= 972891995;
assign addr[12424]= 904098143;
assign addr[12425]= 834157373;
assign addr[12426]= 763158411;
assign addr[12427]= 691191324;
assign addr[12428]= 618347408;
assign addr[12429]= 544719071;
assign addr[12430]= 470399716;
assign addr[12431]= 395483624;
assign addr[12432]= 320065829;
assign addr[12433]= 244242007;
assign addr[12434]= 168108346;
assign addr[12435]= 91761426;
assign addr[12436]= 15298099;
assign addr[12437]= -61184634;
assign addr[12438]= -137589750;
assign addr[12439]= -213820322;
assign addr[12440]= -289779648;
assign addr[12441]= -365371365;
assign addr[12442]= -440499581;
assign addr[12443]= -515068990;
assign addr[12444]= -588984994;
assign addr[12445]= -662153826;
assign addr[12446]= -734482665;
assign addr[12447]= -805879757;
assign addr[12448]= -876254528;
assign addr[12449]= -945517704;
assign addr[12450]= -1013581418;
assign addr[12451]= -1080359326;
assign addr[12452]= -1145766716;
assign addr[12453]= -1209720613;
assign addr[12454]= -1272139887;
assign addr[12455]= -1332945355;
assign addr[12456]= -1392059879;
assign addr[12457]= -1449408469;
assign addr[12458]= -1504918373;
assign addr[12459]= -1558519173;
assign addr[12460]= -1610142873;
assign addr[12461]= -1659723983;
assign addr[12462]= -1707199606;
assign addr[12463]= -1752509516;
assign addr[12464]= -1795596234;
assign addr[12465]= -1836405100;
assign addr[12466]= -1874884346;
assign addr[12467]= -1910985158;
assign addr[12468]= -1944661739;
assign addr[12469]= -1975871368;
assign addr[12470]= -2004574453;
assign addr[12471]= -2030734582;
assign addr[12472]= -2054318569;
assign addr[12473]= -2075296495;
assign addr[12474]= -2093641749;
assign addr[12475]= -2109331059;
assign addr[12476]= -2122344521;
assign addr[12477]= -2132665626;
assign addr[12478]= -2140281282;
assign addr[12479]= -2145181827;
assign addr[12480]= -2147361045;
assign addr[12481]= -2146816171;
assign addr[12482]= -2143547897;
assign addr[12483]= -2137560369;
assign addr[12484]= -2128861181;
assign addr[12485]= -2117461370;
assign addr[12486]= -2103375398;
assign addr[12487]= -2086621133;
assign addr[12488]= -2067219829;
assign addr[12489]= -2045196100;
assign addr[12490]= -2020577882;
assign addr[12491]= -1993396407;
assign addr[12492]= -1963686155;
assign addr[12493]= -1931484818;
assign addr[12494]= -1896833245;
assign addr[12495]= -1859775393;
assign addr[12496]= -1820358275;
assign addr[12497]= -1778631892;
assign addr[12498]= -1734649179;
assign addr[12499]= -1688465931;
assign addr[12500]= -1640140734;
assign addr[12501]= -1589734894;
assign addr[12502]= -1537312353;
assign addr[12503]= -1482939614;
assign addr[12504]= -1426685652;
assign addr[12505]= -1368621831;
assign addr[12506]= -1308821808;
assign addr[12507]= -1247361445;
assign addr[12508]= -1184318708;
assign addr[12509]= -1119773573;
assign addr[12510]= -1053807919;
assign addr[12511]= -986505429;
assign addr[12512]= -917951481;
assign addr[12513]= -848233042;
assign addr[12514]= -777438554;
assign addr[12515]= -705657826;
assign addr[12516]= -632981917;
assign addr[12517]= -559503022;
assign addr[12518]= -485314355;
assign addr[12519]= -410510029;
assign addr[12520]= -335184940;
assign addr[12521]= -259434643;
assign addr[12522]= -183355234;
assign addr[12523]= -107043224;
assign addr[12524]= -30595422;
assign addr[12525]= 45891193;
assign addr[12526]= 122319591;
assign addr[12527]= 198592817;
assign addr[12528]= 274614114;
assign addr[12529]= 350287041;
assign addr[12530]= 425515602;
assign addr[12531]= 500204365;
assign addr[12532]= 574258580;
assign addr[12533]= 647584304;
assign addr[12534]= 720088517;
assign addr[12535]= 791679244;
assign addr[12536]= 862265664;
assign addr[12537]= 931758235;
assign addr[12538]= 1000068799;
assign addr[12539]= 1067110699;
assign addr[12540]= 1132798888;
assign addr[12541]= 1197050035;
assign addr[12542]= 1259782632;
assign addr[12543]= 1320917099;
assign addr[12544]= 1380375881;
assign addr[12545]= 1438083551;
assign addr[12546]= 1493966902;
assign addr[12547]= 1547955041;
assign addr[12548]= 1599979481;
assign addr[12549]= 1649974225;
assign addr[12550]= 1697875851;
assign addr[12551]= 1743623590;
assign addr[12552]= 1787159411;
assign addr[12553]= 1828428082;
assign addr[12554]= 1867377253;
assign addr[12555]= 1903957513;
assign addr[12556]= 1938122457;
assign addr[12557]= 1969828744;
assign addr[12558]= 1999036154;
assign addr[12559]= 2025707632;
assign addr[12560]= 2049809346;
assign addr[12561]= 2071310720;
assign addr[12562]= 2090184478;
assign addr[12563]= 2106406677;
assign addr[12564]= 2119956737;
assign addr[12565]= 2130817471;
assign addr[12566]= 2138975100;
assign addr[12567]= 2144419275;
assign addr[12568]= 2147143090;
assign addr[12569]= 2147143090;
assign addr[12570]= 2144419275;
assign addr[12571]= 2138975100;
assign addr[12572]= 2130817471;
assign addr[12573]= 2119956737;
assign addr[12574]= 2106406677;
assign addr[12575]= 2090184478;
assign addr[12576]= 2071310720;
assign addr[12577]= 2049809346;
assign addr[12578]= 2025707632;
assign addr[12579]= 1999036154;
assign addr[12580]= 1969828744;
assign addr[12581]= 1938122457;
assign addr[12582]= 1903957513;
assign addr[12583]= 1867377253;
assign addr[12584]= 1828428082;
assign addr[12585]= 1787159411;
assign addr[12586]= 1743623590;
assign addr[12587]= 1697875851;
assign addr[12588]= 1649974225;
assign addr[12589]= 1599979481;
assign addr[12590]= 1547955041;
assign addr[12591]= 1493966902;
assign addr[12592]= 1438083551;
assign addr[12593]= 1380375881;
assign addr[12594]= 1320917099;
assign addr[12595]= 1259782632;
assign addr[12596]= 1197050035;
assign addr[12597]= 1132798888;
assign addr[12598]= 1067110699;
assign addr[12599]= 1000068799;
assign addr[12600]= 931758235;
assign addr[12601]= 862265664;
assign addr[12602]= 791679244;
assign addr[12603]= 720088517;
assign addr[12604]= 647584304;
assign addr[12605]= 574258580;
assign addr[12606]= 500204365;
assign addr[12607]= 425515602;
assign addr[12608]= 350287041;
assign addr[12609]= 274614114;
assign addr[12610]= 198592817;
assign addr[12611]= 122319591;
assign addr[12612]= 45891193;
assign addr[12613]= -30595422;
assign addr[12614]= -107043224;
assign addr[12615]= -183355234;
assign addr[12616]= -259434643;
assign addr[12617]= -335184940;
assign addr[12618]= -410510029;
assign addr[12619]= -485314355;
assign addr[12620]= -559503022;
assign addr[12621]= -632981917;
assign addr[12622]= -705657826;
assign addr[12623]= -777438554;
assign addr[12624]= -848233042;
assign addr[12625]= -917951481;
assign addr[12626]= -986505429;
assign addr[12627]= -1053807919;
assign addr[12628]= -1119773573;
assign addr[12629]= -1184318708;
assign addr[12630]= -1247361445;
assign addr[12631]= -1308821808;
assign addr[12632]= -1368621831;
assign addr[12633]= -1426685652;
assign addr[12634]= -1482939614;
assign addr[12635]= -1537312353;
assign addr[12636]= -1589734894;
assign addr[12637]= -1640140734;
assign addr[12638]= -1688465931;
assign addr[12639]= -1734649179;
assign addr[12640]= -1778631892;
assign addr[12641]= -1820358275;
assign addr[12642]= -1859775393;
assign addr[12643]= -1896833245;
assign addr[12644]= -1931484818;
assign addr[12645]= -1963686155;
assign addr[12646]= -1993396407;
assign addr[12647]= -2020577882;
assign addr[12648]= -2045196100;
assign addr[12649]= -2067219829;
assign addr[12650]= -2086621133;
assign addr[12651]= -2103375398;
assign addr[12652]= -2117461370;
assign addr[12653]= -2128861181;
assign addr[12654]= -2137560369;
assign addr[12655]= -2143547897;
assign addr[12656]= -2146816171;
assign addr[12657]= -2147361045;
assign addr[12658]= -2145181827;
assign addr[12659]= -2140281282;
assign addr[12660]= -2132665626;
assign addr[12661]= -2122344521;
assign addr[12662]= -2109331059;
assign addr[12663]= -2093641749;
assign addr[12664]= -2075296495;
assign addr[12665]= -2054318569;
assign addr[12666]= -2030734582;
assign addr[12667]= -2004574453;
assign addr[12668]= -1975871368;
assign addr[12669]= -1944661739;
assign addr[12670]= -1910985158;
assign addr[12671]= -1874884346;
assign addr[12672]= -1836405100;
assign addr[12673]= -1795596234;
assign addr[12674]= -1752509516;
assign addr[12675]= -1707199606;
assign addr[12676]= -1659723983;
assign addr[12677]= -1610142873;
assign addr[12678]= -1558519173;
assign addr[12679]= -1504918373;
assign addr[12680]= -1449408469;
assign addr[12681]= -1392059879;
assign addr[12682]= -1332945355;
assign addr[12683]= -1272139887;
assign addr[12684]= -1209720613;
assign addr[12685]= -1145766716;
assign addr[12686]= -1080359326;
assign addr[12687]= -1013581418;
assign addr[12688]= -945517704;
assign addr[12689]= -876254528;
assign addr[12690]= -805879757;
assign addr[12691]= -734482665;
assign addr[12692]= -662153826;
assign addr[12693]= -588984994;
assign addr[12694]= -515068990;
assign addr[12695]= -440499581;
assign addr[12696]= -365371365;
assign addr[12697]= -289779648;
assign addr[12698]= -213820322;
assign addr[12699]= -137589750;
assign addr[12700]= -61184634;
assign addr[12701]= 15298099;
assign addr[12702]= 91761426;
assign addr[12703]= 168108346;
assign addr[12704]= 244242007;
assign addr[12705]= 320065829;
assign addr[12706]= 395483624;
assign addr[12707]= 470399716;
assign addr[12708]= 544719071;
assign addr[12709]= 618347408;
assign addr[12710]= 691191324;
assign addr[12711]= 763158411;
assign addr[12712]= 834157373;
assign addr[12713]= 904098143;
assign addr[12714]= 972891995;
assign addr[12715]= 1040451659;
assign addr[12716]= 1106691431;
assign addr[12717]= 1171527280;
assign addr[12718]= 1234876957;
assign addr[12719]= 1296660098;
assign addr[12720]= 1356798326;
assign addr[12721]= 1415215352;
assign addr[12722]= 1471837070;
assign addr[12723]= 1526591649;
assign addr[12724]= 1579409630;
assign addr[12725]= 1630224009;
assign addr[12726]= 1678970324;
assign addr[12727]= 1725586737;
assign addr[12728]= 1770014111;
assign addr[12729]= 1812196087;
assign addr[12730]= 1852079154;
assign addr[12731]= 1889612716;
assign addr[12732]= 1924749160;
assign addr[12733]= 1957443913;
assign addr[12734]= 1987655498;
assign addr[12735]= 2015345591;
assign addr[12736]= 2040479063;
assign addr[12737]= 2063024031;
assign addr[12738]= 2082951896;
assign addr[12739]= 2100237377;
assign addr[12740]= 2114858546;
assign addr[12741]= 2126796855;
assign addr[12742]= 2136037160;
assign addr[12743]= 2142567738;
assign addr[12744]= 2146380306;
assign addr[12745]= 2147470025;
assign addr[12746]= 2145835515;
assign addr[12747]= 2141478848;
assign addr[12748]= 2134405552;
assign addr[12749]= 2124624598;
assign addr[12750]= 2112148396;
assign addr[12751]= 2096992772;
assign addr[12752]= 2079176953;
assign addr[12753]= 2058723538;
assign addr[12754]= 2035658475;
assign addr[12755]= 2010011024;
assign addr[12756]= 1981813720;
assign addr[12757]= 1951102334;
assign addr[12758]= 1917915825;
assign addr[12759]= 1882296293;
assign addr[12760]= 1844288924;
assign addr[12761]= 1803941934;
assign addr[12762]= 1761306505;
assign addr[12763]= 1716436725;
assign addr[12764]= 1669389513;
assign addr[12765]= 1620224553;
assign addr[12766]= 1569004214;
assign addr[12767]= 1515793473;
assign addr[12768]= 1460659832;
assign addr[12769]= 1403673233;
assign addr[12770]= 1344905966;
assign addr[12771]= 1284432584;
assign addr[12772]= 1222329801;
assign addr[12773]= 1158676398;
assign addr[12774]= 1093553126;
assign addr[12775]= 1027042599;
assign addr[12776]= 959229189;
assign addr[12777]= 890198924;
assign addr[12778]= 820039373;
assign addr[12779]= 748839539;
assign addr[12780]= 676689746;
assign addr[12781]= 603681519;
assign addr[12782]= 529907477;
assign addr[12783]= 455461206;
assign addr[12784]= 380437148;
assign addr[12785]= 304930476;
assign addr[12786]= 229036977;
assign addr[12787]= 152852926;
assign addr[12788]= 76474970;
assign addr[12789]= 0;
assign addr[12790]= -76474970;
assign addr[12791]= -152852926;
assign addr[12792]= -229036977;
assign addr[12793]= -304930476;
assign addr[12794]= -380437148;
assign addr[12795]= -455461206;
assign addr[12796]= -529907477;
assign addr[12797]= -603681519;
assign addr[12798]= -676689746;
assign addr[12799]= -748839539;
assign addr[12800]= -820039373;
assign addr[12801]= -890198924;
assign addr[12802]= -959229189;
assign addr[12803]= -1027042599;
assign addr[12804]= -1093553126;
assign addr[12805]= -1158676398;
assign addr[12806]= -1222329801;
assign addr[12807]= -1284432584;
assign addr[12808]= -1344905966;
assign addr[12809]= -1403673233;
assign addr[12810]= -1460659832;
assign addr[12811]= -1515793473;
assign addr[12812]= -1569004214;
assign addr[12813]= -1620224553;
assign addr[12814]= -1669389513;
assign addr[12815]= -1716436725;
assign addr[12816]= -1761306505;
assign addr[12817]= -1803941934;
assign addr[12818]= -1844288924;
assign addr[12819]= -1882296293;
assign addr[12820]= -1917915825;
assign addr[12821]= -1951102334;
assign addr[12822]= -1981813720;
assign addr[12823]= -2010011024;
assign addr[12824]= -2035658475;
assign addr[12825]= -2058723538;
assign addr[12826]= -2079176953;
assign addr[12827]= -2096992772;
assign addr[12828]= -2112148396;
assign addr[12829]= -2124624598;
assign addr[12830]= -2134405552;
assign addr[12831]= -2141478848;
assign addr[12832]= -2145835515;
assign addr[12833]= -2147470025;
assign addr[12834]= -2146380306;
assign addr[12835]= -2142567738;
assign addr[12836]= -2136037160;
assign addr[12837]= -2126796855;
assign addr[12838]= -2114858546;
assign addr[12839]= -2100237377;
assign addr[12840]= -2082951896;
assign addr[12841]= -2063024031;
assign addr[12842]= -2040479063;
assign addr[12843]= -2015345591;
assign addr[12844]= -1987655498;
assign addr[12845]= -1957443913;
assign addr[12846]= -1924749160;
assign addr[12847]= -1889612716;
assign addr[12848]= -1852079154;
assign addr[12849]= -1812196087;
assign addr[12850]= -1770014111;
assign addr[12851]= -1725586737;
assign addr[12852]= -1678970324;
assign addr[12853]= -1630224009;
assign addr[12854]= -1579409630;
assign addr[12855]= -1526591649;
assign addr[12856]= -1471837070;
assign addr[12857]= -1415215352;
assign addr[12858]= -1356798326;
assign addr[12859]= -1296660098;
assign addr[12860]= -1234876957;
assign addr[12861]= -1171527280;
assign addr[12862]= -1106691431;
assign addr[12863]= -1040451659;
assign addr[12864]= -972891995;
assign addr[12865]= -904098143;
assign addr[12866]= -834157373;
assign addr[12867]= -763158411;
assign addr[12868]= -691191324;
assign addr[12869]= -618347408;
assign addr[12870]= -544719071;
assign addr[12871]= -470399716;
assign addr[12872]= -395483624;
assign addr[12873]= -320065829;
assign addr[12874]= -244242007;
assign addr[12875]= -168108346;
assign addr[12876]= -91761426;
assign addr[12877]= -15298099;
assign addr[12878]= 61184634;
assign addr[12879]= 137589750;
assign addr[12880]= 213820322;
assign addr[12881]= 289779648;
assign addr[12882]= 365371365;
assign addr[12883]= 440499581;
assign addr[12884]= 515068990;
assign addr[12885]= 588984994;
assign addr[12886]= 662153826;
assign addr[12887]= 734482665;
assign addr[12888]= 805879757;
assign addr[12889]= 876254528;
assign addr[12890]= 945517704;
assign addr[12891]= 1013581418;
assign addr[12892]= 1080359326;
assign addr[12893]= 1145766716;
assign addr[12894]= 1209720613;
assign addr[12895]= 1272139887;
assign addr[12896]= 1332945355;
assign addr[12897]= 1392059879;
assign addr[12898]= 1449408469;
assign addr[12899]= 1504918373;
assign addr[12900]= 1558519173;
assign addr[12901]= 1610142873;
assign addr[12902]= 1659723983;
assign addr[12903]= 1707199606;
assign addr[12904]= 1752509516;
assign addr[12905]= 1795596234;
assign addr[12906]= 1836405100;
assign addr[12907]= 1874884346;
assign addr[12908]= 1910985158;
assign addr[12909]= 1944661739;
assign addr[12910]= 1975871368;
assign addr[12911]= 2004574453;
assign addr[12912]= 2030734582;
assign addr[12913]= 2054318569;
assign addr[12914]= 2075296495;
assign addr[12915]= 2093641749;
assign addr[12916]= 2109331059;
assign addr[12917]= 2122344521;
assign addr[12918]= 2132665626;
assign addr[12919]= 2140281282;
assign addr[12920]= 2145181827;
assign addr[12921]= 2147361045;
assign addr[12922]= 2146816171;
assign addr[12923]= 2143547897;
assign addr[12924]= 2137560369;
assign addr[12925]= 2128861181;
assign addr[12926]= 2117461370;
assign addr[12927]= 2103375398;
assign addr[12928]= 2086621133;
assign addr[12929]= 2067219829;
assign addr[12930]= 2045196100;
assign addr[12931]= 2020577882;
assign addr[12932]= 1993396407;
assign addr[12933]= 1963686155;
assign addr[12934]= 1931484818;
assign addr[12935]= 1896833245;
assign addr[12936]= 1859775393;
assign addr[12937]= 1820358275;
assign addr[12938]= 1778631892;
assign addr[12939]= 1734649179;
assign addr[12940]= 1688465931;
assign addr[12941]= 1640140734;
assign addr[12942]= 1589734894;
assign addr[12943]= 1537312353;
assign addr[12944]= 1482939614;
assign addr[12945]= 1426685652;
assign addr[12946]= 1368621831;
assign addr[12947]= 1308821808;
assign addr[12948]= 1247361445;
assign addr[12949]= 1184318708;
assign addr[12950]= 1119773573;
assign addr[12951]= 1053807919;
assign addr[12952]= 986505429;
assign addr[12953]= 917951481;
assign addr[12954]= 848233042;
assign addr[12955]= 777438554;
assign addr[12956]= 705657826;
assign addr[12957]= 632981917;
assign addr[12958]= 559503022;
assign addr[12959]= 485314355;
assign addr[12960]= 410510029;
assign addr[12961]= 335184940;
assign addr[12962]= 259434643;
assign addr[12963]= 183355234;
assign addr[12964]= 107043224;
assign addr[12965]= 30595422;
assign addr[12966]= -45891193;
assign addr[12967]= -122319591;
assign addr[12968]= -198592817;
assign addr[12969]= -274614114;
assign addr[12970]= -350287041;
assign addr[12971]= -425515602;
assign addr[12972]= -500204365;
assign addr[12973]= -574258580;
assign addr[12974]= -647584304;
assign addr[12975]= -720088517;
assign addr[12976]= -791679244;
assign addr[12977]= -862265664;
assign addr[12978]= -931758235;
assign addr[12979]= -1000068799;
assign addr[12980]= -1067110699;
assign addr[12981]= -1132798888;
assign addr[12982]= -1197050035;
assign addr[12983]= -1259782632;
assign addr[12984]= -1320917099;
assign addr[12985]= -1380375881;
assign addr[12986]= -1438083551;
assign addr[12987]= -1493966902;
assign addr[12988]= -1547955041;
assign addr[12989]= -1599979481;
assign addr[12990]= -1649974225;
assign addr[12991]= -1697875851;
assign addr[12992]= -1743623590;
assign addr[12993]= -1787159411;
assign addr[12994]= -1828428082;
assign addr[12995]= -1867377253;
assign addr[12996]= -1903957513;
assign addr[12997]= -1938122457;
assign addr[12998]= -1969828744;
assign addr[12999]= -1999036154;
assign addr[13000]= -2025707632;
assign addr[13001]= -2049809346;
assign addr[13002]= -2071310720;
assign addr[13003]= -2090184478;
assign addr[13004]= -2106406677;
assign addr[13005]= -2119956737;
assign addr[13006]= -2130817471;
assign addr[13007]= -2138975100;
assign addr[13008]= -2144419275;
assign addr[13009]= -2147143090;
assign addr[13010]= -2147143090;
assign addr[13011]= -2144419275;
assign addr[13012]= -2138975100;
assign addr[13013]= -2130817471;
assign addr[13014]= -2119956737;
assign addr[13015]= -2106406677;
assign addr[13016]= -2090184478;
assign addr[13017]= -2071310720;
assign addr[13018]= -2049809346;
assign addr[13019]= -2025707632;
assign addr[13020]= -1999036154;
assign addr[13021]= -1969828744;
assign addr[13022]= -1938122457;
assign addr[13023]= -1903957513;
assign addr[13024]= -1867377253;
assign addr[13025]= -1828428082;
assign addr[13026]= -1787159411;
assign addr[13027]= -1743623590;
assign addr[13028]= -1697875851;
assign addr[13029]= -1649974225;
assign addr[13030]= -1599979481;
assign addr[13031]= -1547955041;
assign addr[13032]= -1493966902;
assign addr[13033]= -1438083551;
assign addr[13034]= -1380375881;
assign addr[13035]= -1320917099;
assign addr[13036]= -1259782632;
assign addr[13037]= -1197050035;
assign addr[13038]= -1132798888;
assign addr[13039]= -1067110699;
assign addr[13040]= -1000068799;
assign addr[13041]= -931758235;
assign addr[13042]= -862265664;
assign addr[13043]= -791679244;
assign addr[13044]= -720088517;
assign addr[13045]= -647584304;
assign addr[13046]= -574258580;
assign addr[13047]= -500204365;
assign addr[13048]= -425515602;
assign addr[13049]= -350287041;
assign addr[13050]= -274614114;
assign addr[13051]= -198592817;
assign addr[13052]= -122319591;
assign addr[13053]= -45891193;
assign addr[13054]= 30595422;
assign addr[13055]= 107043224;
assign addr[13056]= 183355234;
assign addr[13057]= 259434643;
assign addr[13058]= 335184940;
assign addr[13059]= 410510029;
assign addr[13060]= 485314355;
assign addr[13061]= 559503022;
assign addr[13062]= 632981917;
assign addr[13063]= 705657826;
assign addr[13064]= 777438554;
assign addr[13065]= 848233042;
assign addr[13066]= 917951481;
assign addr[13067]= 986505429;
assign addr[13068]= 1053807919;
assign addr[13069]= 1119773573;
assign addr[13070]= 1184318708;
assign addr[13071]= 1247361445;
assign addr[13072]= 1308821808;
assign addr[13073]= 1368621831;
assign addr[13074]= 1426685652;
assign addr[13075]= 1482939614;
assign addr[13076]= 1537312353;
assign addr[13077]= 1589734894;
assign addr[13078]= 1640140734;
assign addr[13079]= 1688465931;
assign addr[13080]= 1734649179;
assign addr[13081]= 1778631892;
assign addr[13082]= 1820358275;
assign addr[13083]= 1859775393;
assign addr[13084]= 1896833245;
assign addr[13085]= 1931484818;
assign addr[13086]= 1963686155;
assign addr[13087]= 1993396407;
assign addr[13088]= 2020577882;
assign addr[13089]= 2045196100;
assign addr[13090]= 2067219829;
assign addr[13091]= 2086621133;
assign addr[13092]= 2103375398;
assign addr[13093]= 2117461370;
assign addr[13094]= 2128861181;
assign addr[13095]= 2137560369;
assign addr[13096]= 2143547897;
assign addr[13097]= 2146816171;
assign addr[13098]= 2147361045;
assign addr[13099]= 2145181827;
assign addr[13100]= 2140281282;
assign addr[13101]= 2132665626;
assign addr[13102]= 2122344521;
assign addr[13103]= 2109331059;
assign addr[13104]= 2093641749;
assign addr[13105]= 2075296495;
assign addr[13106]= 2054318569;
assign addr[13107]= 2030734582;
assign addr[13108]= 2004574453;
assign addr[13109]= 1975871368;
assign addr[13110]= 1944661739;
assign addr[13111]= 1910985158;
assign addr[13112]= 1874884346;
assign addr[13113]= 1836405100;
assign addr[13114]= 1795596234;
assign addr[13115]= 1752509516;
assign addr[13116]= 1707199606;
assign addr[13117]= 1659723983;
assign addr[13118]= 1610142873;
assign addr[13119]= 1558519173;
assign addr[13120]= 1504918373;
assign addr[13121]= 1449408469;
assign addr[13122]= 1392059879;
assign addr[13123]= 1332945355;
assign addr[13124]= 1272139887;
assign addr[13125]= 1209720613;
assign addr[13126]= 1145766716;
assign addr[13127]= 1080359326;
assign addr[13128]= 1013581418;
assign addr[13129]= 945517704;
assign addr[13130]= 876254528;
assign addr[13131]= 805879757;
assign addr[13132]= 734482665;
assign addr[13133]= 662153826;
assign addr[13134]= 588984994;
assign addr[13135]= 515068990;
assign addr[13136]= 440499581;
assign addr[13137]= 365371365;
assign addr[13138]= 289779648;
assign addr[13139]= 213820322;
assign addr[13140]= 137589750;
assign addr[13141]= 61184634;
assign addr[13142]= -15298099;
assign addr[13143]= -91761426;
assign addr[13144]= -168108346;
assign addr[13145]= -244242007;
assign addr[13146]= -320065829;
assign addr[13147]= -395483624;
assign addr[13148]= -470399716;
assign addr[13149]= -544719071;
assign addr[13150]= -618347408;
assign addr[13151]= -691191324;
assign addr[13152]= -763158411;
assign addr[13153]= -834157373;
assign addr[13154]= -904098143;
assign addr[13155]= -972891995;
assign addr[13156]= -1040451659;
assign addr[13157]= -1106691431;
assign addr[13158]= -1171527280;
assign addr[13159]= -1234876957;
assign addr[13160]= -1296660098;
assign addr[13161]= -1356798326;
assign addr[13162]= -1415215352;
assign addr[13163]= -1471837070;
assign addr[13164]= -1526591649;
assign addr[13165]= -1579409630;
assign addr[13166]= -1630224009;
assign addr[13167]= -1678970324;
assign addr[13168]= -1725586737;
assign addr[13169]= -1770014111;
assign addr[13170]= -1812196087;
assign addr[13171]= -1852079154;
assign addr[13172]= -1889612716;
assign addr[13173]= -1924749160;
assign addr[13174]= -1957443913;
assign addr[13175]= -1987655498;
assign addr[13176]= -2015345591;
assign addr[13177]= -2040479063;
assign addr[13178]= -2063024031;
assign addr[13179]= -2082951896;
assign addr[13180]= -2100237377;
assign addr[13181]= -2114858546;
assign addr[13182]= -2126796855;
assign addr[13183]= -2136037160;
assign addr[13184]= -2142567738;
assign addr[13185]= -2146380306;
assign addr[13186]= -2147470025;
assign addr[13187]= -2145835515;
assign addr[13188]= -2141478848;
assign addr[13189]= -2134405552;
assign addr[13190]= -2124624598;
assign addr[13191]= -2112148396;
assign addr[13192]= -2096992772;
assign addr[13193]= -2079176953;
assign addr[13194]= -2058723538;
assign addr[13195]= -2035658475;
assign addr[13196]= -2010011024;
assign addr[13197]= -1981813720;
assign addr[13198]= -1951102334;
assign addr[13199]= -1917915825;
assign addr[13200]= -1882296293;
assign addr[13201]= -1844288924;
assign addr[13202]= -1803941934;
assign addr[13203]= -1761306505;
assign addr[13204]= -1716436725;
assign addr[13205]= -1669389513;
assign addr[13206]= -1620224553;
assign addr[13207]= -1569004214;
assign addr[13208]= -1515793473;
assign addr[13209]= -1460659832;
assign addr[13210]= -1403673233;
assign addr[13211]= -1344905966;
assign addr[13212]= -1284432584;
assign addr[13213]= -1222329801;
assign addr[13214]= -1158676398;
assign addr[13215]= -1093553126;
assign addr[13216]= -1027042599;
assign addr[13217]= -959229189;
assign addr[13218]= -890198924;
assign addr[13219]= -820039373;
assign addr[13220]= -748839539;
assign addr[13221]= -676689746;
assign addr[13222]= -603681519;
assign addr[13223]= -529907477;
assign addr[13224]= -455461206;
assign addr[13225]= -380437148;
assign addr[13226]= -304930476;
assign addr[13227]= -229036977;
assign addr[13228]= -152852926;
assign addr[13229]= -76474970;
assign addr[13230]= 0;
assign addr[13231]= 76474970;
assign addr[13232]= 152852926;
assign addr[13233]= 229036977;
assign addr[13234]= 304930476;
assign addr[13235]= 380437148;
assign addr[13236]= 455461206;
assign addr[13237]= 529907477;
assign addr[13238]= 603681519;
assign addr[13239]= 676689746;
assign addr[13240]= 748839539;
assign addr[13241]= 820039373;
assign addr[13242]= 890198924;
assign addr[13243]= 959229189;
assign addr[13244]= 1027042599;
assign addr[13245]= 1093553126;
assign addr[13246]= 1158676398;
assign addr[13247]= 1222329801;
assign addr[13248]= 1284432584;
assign addr[13249]= 1344905966;
assign addr[13250]= 1403673233;
assign addr[13251]= 1460659832;
assign addr[13252]= 1515793473;
assign addr[13253]= 1569004214;
assign addr[13254]= 1620224553;
assign addr[13255]= 1669389513;
assign addr[13256]= 1716436725;
assign addr[13257]= 1761306505;
assign addr[13258]= 1803941934;
assign addr[13259]= 1844288924;
assign addr[13260]= 1882296293;
assign addr[13261]= 1917915825;
assign addr[13262]= 1951102334;
assign addr[13263]= 1981813720;
assign addr[13264]= 2010011024;
assign addr[13265]= 2035658475;
assign addr[13266]= 2058723538;
assign addr[13267]= 2079176953;
assign addr[13268]= 2096992772;
assign addr[13269]= 2112148396;
assign addr[13270]= 2124624598;
assign addr[13271]= 2134405552;
assign addr[13272]= 2141478848;
assign addr[13273]= 2145835515;
assign addr[13274]= 2147470025;
assign addr[13275]= 2146380306;
assign addr[13276]= 2142567738;
assign addr[13277]= 2136037160;
assign addr[13278]= 2126796855;
assign addr[13279]= 2114858546;
assign addr[13280]= 2100237377;
assign addr[13281]= 2082951896;
assign addr[13282]= 2063024031;
assign addr[13283]= 2040479063;
assign addr[13284]= 2015345591;
assign addr[13285]= 1987655498;
assign addr[13286]= 1957443913;
assign addr[13287]= 1924749160;
assign addr[13288]= 1889612716;
assign addr[13289]= 1852079154;
assign addr[13290]= 1812196087;
assign addr[13291]= 1770014111;
assign addr[13292]= 1725586737;
assign addr[13293]= 1678970324;
assign addr[13294]= 1630224009;
assign addr[13295]= 1579409630;
assign addr[13296]= 1526591649;
assign addr[13297]= 1471837070;
assign addr[13298]= 1415215352;
assign addr[13299]= 1356798326;
assign addr[13300]= 1296660098;
assign addr[13301]= 1234876957;
assign addr[13302]= 1171527280;
assign addr[13303]= 1106691431;
assign addr[13304]= 1040451659;
assign addr[13305]= 972891995;
assign addr[13306]= 904098143;
assign addr[13307]= 834157373;
assign addr[13308]= 763158411;
assign addr[13309]= 691191324;
assign addr[13310]= 618347408;
assign addr[13311]= 544719071;
assign addr[13312]= 470399716;
assign addr[13313]= 395483624;
assign addr[13314]= 320065829;
assign addr[13315]= 244242007;
assign addr[13316]= 168108346;
assign addr[13317]= 91761426;
assign addr[13318]= 15298099;
assign addr[13319]= -61184634;
assign addr[13320]= -137589750;
assign addr[13321]= -213820322;
assign addr[13322]= -289779648;
assign addr[13323]= -365371365;
assign addr[13324]= -440499581;
assign addr[13325]= -515068990;
assign addr[13326]= -588984994;
assign addr[13327]= -662153826;
assign addr[13328]= -734482665;
assign addr[13329]= -805879757;
assign addr[13330]= -876254528;
assign addr[13331]= -945517704;
assign addr[13332]= -1013581418;
assign addr[13333]= -1080359326;
assign addr[13334]= -1145766716;
assign addr[13335]= -1209720613;
assign addr[13336]= -1272139887;
assign addr[13337]= -1332945355;
assign addr[13338]= -1392059879;
assign addr[13339]= -1449408469;
assign addr[13340]= -1504918373;
assign addr[13341]= -1558519173;
assign addr[13342]= -1610142873;
assign addr[13343]= -1659723983;
assign addr[13344]= -1707199606;
assign addr[13345]= -1752509516;
assign addr[13346]= -1795596234;
assign addr[13347]= -1836405100;
assign addr[13348]= -1874884346;
assign addr[13349]= -1910985158;
assign addr[13350]= -1944661739;
assign addr[13351]= -1975871368;
assign addr[13352]= -2004574453;
assign addr[13353]= -2030734582;
assign addr[13354]= -2054318569;
assign addr[13355]= -2075296495;
assign addr[13356]= -2093641749;
assign addr[13357]= -2109331059;
assign addr[13358]= -2122344521;
assign addr[13359]= -2132665626;
assign addr[13360]= -2140281282;
assign addr[13361]= -2145181827;
assign addr[13362]= -2147361045;
assign addr[13363]= -2146816171;
assign addr[13364]= -2143547897;
assign addr[13365]= -2137560369;
assign addr[13366]= -2128861181;
assign addr[13367]= -2117461370;
assign addr[13368]= -2103375398;
assign addr[13369]= -2086621133;
assign addr[13370]= -2067219829;
assign addr[13371]= -2045196100;
assign addr[13372]= -2020577882;
assign addr[13373]= -1993396407;
assign addr[13374]= -1963686155;
assign addr[13375]= -1931484818;
assign addr[13376]= -1896833245;
assign addr[13377]= -1859775393;
assign addr[13378]= -1820358275;
assign addr[13379]= -1778631892;
assign addr[13380]= -1734649179;
assign addr[13381]= -1688465931;
assign addr[13382]= -1640140734;
assign addr[13383]= -1589734894;
assign addr[13384]= -1537312353;
assign addr[13385]= -1482939614;
assign addr[13386]= -1426685652;
assign addr[13387]= -1368621831;
assign addr[13388]= -1308821808;
assign addr[13389]= -1247361445;
assign addr[13390]= -1184318708;
assign addr[13391]= -1119773573;
assign addr[13392]= -1053807919;
assign addr[13393]= -986505429;
assign addr[13394]= -917951481;
assign addr[13395]= -848233042;
assign addr[13396]= -777438554;
assign addr[13397]= -705657826;
assign addr[13398]= -632981917;
assign addr[13399]= -559503022;
assign addr[13400]= -485314355;
assign addr[13401]= -410510029;
assign addr[13402]= -335184940;
assign addr[13403]= -259434643;
assign addr[13404]= -183355234;
assign addr[13405]= -107043224;
assign addr[13406]= -30595422;
assign addr[13407]= 45891193;
assign addr[13408]= 122319591;
assign addr[13409]= 198592817;
assign addr[13410]= 274614114;
assign addr[13411]= 350287041;
assign addr[13412]= 425515602;
assign addr[13413]= 500204365;
assign addr[13414]= 574258580;
assign addr[13415]= 647584304;
assign addr[13416]= 720088517;
assign addr[13417]= 791679244;
assign addr[13418]= 862265664;
assign addr[13419]= 931758235;
assign addr[13420]= 1000068799;
assign addr[13421]= 1067110699;
assign addr[13422]= 1132798888;
assign addr[13423]= 1197050035;
assign addr[13424]= 1259782632;
assign addr[13425]= 1320917099;
assign addr[13426]= 1380375881;
assign addr[13427]= 1438083551;
assign addr[13428]= 1493966902;
assign addr[13429]= 1547955041;
assign addr[13430]= 1599979481;
assign addr[13431]= 1649974225;
assign addr[13432]= 1697875851;
assign addr[13433]= 1743623590;
assign addr[13434]= 1787159411;
assign addr[13435]= 1828428082;
assign addr[13436]= 1867377253;
assign addr[13437]= 1903957513;
assign addr[13438]= 1938122457;
assign addr[13439]= 1969828744;
assign addr[13440]= 1999036154;
assign addr[13441]= 2025707632;
assign addr[13442]= 2049809346;
assign addr[13443]= 2071310720;
assign addr[13444]= 2090184478;
assign addr[13445]= 2106406677;
assign addr[13446]= 2119956737;
assign addr[13447]= 2130817471;
assign addr[13448]= 2138975100;
assign addr[13449]= 2144419275;
assign addr[13450]= 2147143090;
assign addr[13451]= 2147143090;
assign addr[13452]= 2144419275;
assign addr[13453]= 2138975100;
assign addr[13454]= 2130817471;
assign addr[13455]= 2119956737;
assign addr[13456]= 2106406677;
assign addr[13457]= 2090184478;
assign addr[13458]= 2071310720;
assign addr[13459]= 2049809346;
assign addr[13460]= 2025707632;
assign addr[13461]= 1999036154;
assign addr[13462]= 1969828744;
assign addr[13463]= 1938122457;
assign addr[13464]= 1903957513;
assign addr[13465]= 1867377253;
assign addr[13466]= 1828428082;
assign addr[13467]= 1787159411;
assign addr[13468]= 1743623590;
assign addr[13469]= 1697875851;
assign addr[13470]= 1649974225;
assign addr[13471]= 1599979481;
assign addr[13472]= 1547955041;
assign addr[13473]= 1493966902;
assign addr[13474]= 1438083551;
assign addr[13475]= 1380375881;
assign addr[13476]= 1320917099;
assign addr[13477]= 1259782632;
assign addr[13478]= 1197050035;
assign addr[13479]= 1132798888;
assign addr[13480]= 1067110699;
assign addr[13481]= 1000068799;
assign addr[13482]= 931758235;
assign addr[13483]= 862265664;
assign addr[13484]= 791679244;
assign addr[13485]= 720088517;
assign addr[13486]= 647584304;
assign addr[13487]= 574258580;
assign addr[13488]= 500204365;
assign addr[13489]= 425515602;
assign addr[13490]= 350287041;
assign addr[13491]= 274614114;
assign addr[13492]= 198592817;
assign addr[13493]= 122319591;
assign addr[13494]= 45891193;
assign addr[13495]= -30595422;
assign addr[13496]= -107043224;
assign addr[13497]= -183355234;
assign addr[13498]= -259434643;
assign addr[13499]= -335184940;
assign addr[13500]= -410510029;
assign addr[13501]= -485314355;
assign addr[13502]= -559503022;
assign addr[13503]= -632981917;
assign addr[13504]= -705657826;
assign addr[13505]= -777438554;
assign addr[13506]= -848233042;
assign addr[13507]= -917951481;
assign addr[13508]= -986505429;
assign addr[13509]= -1053807919;
assign addr[13510]= -1119773573;
assign addr[13511]= -1184318708;
assign addr[13512]= -1247361445;
assign addr[13513]= -1308821808;
assign addr[13514]= -1368621831;
assign addr[13515]= -1426685652;
assign addr[13516]= -1482939614;
assign addr[13517]= -1537312353;
assign addr[13518]= -1589734894;
assign addr[13519]= -1640140734;
assign addr[13520]= -1688465931;
assign addr[13521]= -1734649179;
assign addr[13522]= -1778631892;
assign addr[13523]= -1820358275;
assign addr[13524]= -1859775393;
assign addr[13525]= -1896833245;
assign addr[13526]= -1931484818;
assign addr[13527]= -1963686155;
assign addr[13528]= -1993396407;
assign addr[13529]= -2020577882;
assign addr[13530]= -2045196100;
assign addr[13531]= -2067219829;
assign addr[13532]= -2086621133;
assign addr[13533]= -2103375398;
assign addr[13534]= -2117461370;
assign addr[13535]= -2128861181;
assign addr[13536]= -2137560369;
assign addr[13537]= -2143547897;
assign addr[13538]= -2146816171;
assign addr[13539]= -2147361045;
assign addr[13540]= -2145181827;
assign addr[13541]= -2140281282;
assign addr[13542]= -2132665626;
assign addr[13543]= -2122344521;
assign addr[13544]= -2109331059;
assign addr[13545]= -2093641749;
assign addr[13546]= -2075296495;
assign addr[13547]= -2054318569;
assign addr[13548]= -2030734582;
assign addr[13549]= -2004574453;
assign addr[13550]= -1975871368;
assign addr[13551]= -1944661739;
assign addr[13552]= -1910985158;
assign addr[13553]= -1874884346;
assign addr[13554]= -1836405100;
assign addr[13555]= -1795596234;
assign addr[13556]= -1752509516;
assign addr[13557]= -1707199606;
assign addr[13558]= -1659723983;
assign addr[13559]= -1610142873;
assign addr[13560]= -1558519173;
assign addr[13561]= -1504918373;
assign addr[13562]= -1449408469;
assign addr[13563]= -1392059879;
assign addr[13564]= -1332945355;
assign addr[13565]= -1272139887;
assign addr[13566]= -1209720613;
assign addr[13567]= -1145766716;
assign addr[13568]= -1080359326;
assign addr[13569]= -1013581418;
assign addr[13570]= -945517704;
assign addr[13571]= -876254528;
assign addr[13572]= -805879757;
assign addr[13573]= -734482665;
assign addr[13574]= -662153826;
assign addr[13575]= -588984994;
assign addr[13576]= -515068990;
assign addr[13577]= -440499581;
assign addr[13578]= -365371365;
assign addr[13579]= -289779648;
assign addr[13580]= -213820322;
assign addr[13581]= -137589750;
assign addr[13582]= -61184634;
assign addr[13583]= 15298099;
assign addr[13584]= 91761426;
assign addr[13585]= 168108346;
assign addr[13586]= 244242007;
assign addr[13587]= 320065829;
assign addr[13588]= 395483624;
assign addr[13589]= 470399716;
assign addr[13590]= 544719071;
assign addr[13591]= 618347408;
assign addr[13592]= 691191324;
assign addr[13593]= 763158411;
assign addr[13594]= 834157373;
assign addr[13595]= 904098143;
assign addr[13596]= 972891995;
assign addr[13597]= 1040451659;
assign addr[13598]= 1106691431;
assign addr[13599]= 1171527280;
assign addr[13600]= 1234876957;
assign addr[13601]= 1296660098;
assign addr[13602]= 1356798326;
assign addr[13603]= 1415215352;
assign addr[13604]= 1471837070;
assign addr[13605]= 1526591649;
assign addr[13606]= 1579409630;
assign addr[13607]= 1630224009;
assign addr[13608]= 1678970324;
assign addr[13609]= 1725586737;
assign addr[13610]= 1770014111;
assign addr[13611]= 1812196087;
assign addr[13612]= 1852079154;
assign addr[13613]= 1889612716;
assign addr[13614]= 1924749160;
assign addr[13615]= 1957443913;
assign addr[13616]= 1987655498;
assign addr[13617]= 2015345591;
assign addr[13618]= 2040479063;
assign addr[13619]= 2063024031;
assign addr[13620]= 2082951896;
assign addr[13621]= 2100237377;
assign addr[13622]= 2114858546;
assign addr[13623]= 2126796855;
assign addr[13624]= 2136037160;
assign addr[13625]= 2142567738;
assign addr[13626]= 2146380306;
assign addr[13627]= 2147470025;
assign addr[13628]= 2145835515;
assign addr[13629]= 2141478848;
assign addr[13630]= 2134405552;
assign addr[13631]= 2124624598;
assign addr[13632]= 2112148396;
assign addr[13633]= 2096992772;
assign addr[13634]= 2079176953;
assign addr[13635]= 2058723538;
assign addr[13636]= 2035658475;
assign addr[13637]= 2010011024;
assign addr[13638]= 1981813720;
assign addr[13639]= 1951102334;
assign addr[13640]= 1917915825;
assign addr[13641]= 1882296293;
assign addr[13642]= 1844288924;
assign addr[13643]= 1803941934;
assign addr[13644]= 1761306505;
assign addr[13645]= 1716436725;
assign addr[13646]= 1669389513;
assign addr[13647]= 1620224553;
assign addr[13648]= 1569004214;
assign addr[13649]= 1515793473;
assign addr[13650]= 1460659832;
assign addr[13651]= 1403673233;
assign addr[13652]= 1344905966;
assign addr[13653]= 1284432584;
assign addr[13654]= 1222329801;
assign addr[13655]= 1158676398;
assign addr[13656]= 1093553126;
assign addr[13657]= 1027042599;
assign addr[13658]= 959229189;
assign addr[13659]= 890198924;
assign addr[13660]= 820039373;
assign addr[13661]= 748839539;
assign addr[13662]= 676689746;
assign addr[13663]= 603681519;
assign addr[13664]= 529907477;
assign addr[13665]= 455461206;
assign addr[13666]= 380437148;
assign addr[13667]= 304930476;
assign addr[13668]= 229036977;
assign addr[13669]= 152852926;
assign addr[13670]= 76474970;
assign addr[13671]= 0;
assign addr[13672]= -76474970;
assign addr[13673]= -152852926;
assign addr[13674]= -229036977;
assign addr[13675]= -304930476;
assign addr[13676]= -380437148;
assign addr[13677]= -455461206;
assign addr[13678]= -529907477;
assign addr[13679]= -603681519;
assign addr[13680]= -676689746;
assign addr[13681]= -748839539;
assign addr[13682]= -820039373;
assign addr[13683]= -890198924;
assign addr[13684]= -959229189;
assign addr[13685]= -1027042599;
assign addr[13686]= -1093553126;
assign addr[13687]= -1158676398;
assign addr[13688]= -1222329801;
assign addr[13689]= -1284432584;
assign addr[13690]= -1344905966;
assign addr[13691]= -1403673233;
assign addr[13692]= -1460659832;
assign addr[13693]= -1515793473;
assign addr[13694]= -1569004214;
assign addr[13695]= -1620224553;
assign addr[13696]= -1669389513;
assign addr[13697]= -1716436725;
assign addr[13698]= -1761306505;
assign addr[13699]= -1803941934;
assign addr[13700]= -1844288924;
assign addr[13701]= -1882296293;
assign addr[13702]= -1917915825;
assign addr[13703]= -1951102334;
assign addr[13704]= -1981813720;
assign addr[13705]= -2010011024;
assign addr[13706]= -2035658475;
assign addr[13707]= -2058723538;
assign addr[13708]= -2079176953;
assign addr[13709]= -2096992772;
assign addr[13710]= -2112148396;
assign addr[13711]= -2124624598;
assign addr[13712]= -2134405552;
assign addr[13713]= -2141478848;
assign addr[13714]= -2145835515;
assign addr[13715]= -2147470025;
assign addr[13716]= -2146380306;
assign addr[13717]= -2142567738;
assign addr[13718]= -2136037160;
assign addr[13719]= -2126796855;
assign addr[13720]= -2114858546;
assign addr[13721]= -2100237377;
assign addr[13722]= -2082951896;
assign addr[13723]= -2063024031;
assign addr[13724]= -2040479063;
assign addr[13725]= -2015345591;
assign addr[13726]= -1987655498;
assign addr[13727]= -1957443913;
assign addr[13728]= -1924749160;
assign addr[13729]= -1889612716;
assign addr[13730]= -1852079154;
assign addr[13731]= -1812196087;
assign addr[13732]= -1770014111;
assign addr[13733]= -1725586737;
assign addr[13734]= -1678970324;
assign addr[13735]= -1630224009;
assign addr[13736]= -1579409630;
assign addr[13737]= -1526591649;
assign addr[13738]= -1471837070;
assign addr[13739]= -1415215352;
assign addr[13740]= -1356798326;
assign addr[13741]= -1296660098;
assign addr[13742]= -1234876957;
assign addr[13743]= -1171527280;
assign addr[13744]= -1106691431;
assign addr[13745]= -1040451659;
assign addr[13746]= -972891995;
assign addr[13747]= -904098143;
assign addr[13748]= -834157373;
assign addr[13749]= -763158411;
assign addr[13750]= -691191324;
assign addr[13751]= -618347408;
assign addr[13752]= -544719071;
assign addr[13753]= -470399716;
assign addr[13754]= -395483624;
assign addr[13755]= -320065829;
assign addr[13756]= -244242007;
assign addr[13757]= -168108346;
assign addr[13758]= -91761426;
assign addr[13759]= -15298099;
assign addr[13760]= 61184634;
assign addr[13761]= 137589750;
assign addr[13762]= 213820322;
assign addr[13763]= 289779648;
assign addr[13764]= 365371365;
assign addr[13765]= 440499581;
assign addr[13766]= 515068990;
assign addr[13767]= 588984994;
assign addr[13768]= 662153826;
assign addr[13769]= 734482665;
assign addr[13770]= 805879757;
assign addr[13771]= 876254528;
assign addr[13772]= 945517704;
assign addr[13773]= 1013581418;
assign addr[13774]= 1080359326;
assign addr[13775]= 1145766716;
assign addr[13776]= 1209720613;
assign addr[13777]= 1272139887;
assign addr[13778]= 1332945355;
assign addr[13779]= 1392059879;
assign addr[13780]= 1449408469;
assign addr[13781]= 1504918373;
assign addr[13782]= 1558519173;
assign addr[13783]= 1610142873;
assign addr[13784]= 1659723983;
assign addr[13785]= 1707199606;
assign addr[13786]= 1752509516;
assign addr[13787]= 1795596234;
assign addr[13788]= 1836405100;
assign addr[13789]= 1874884346;
assign addr[13790]= 1910985158;
assign addr[13791]= 1944661739;
assign addr[13792]= 1975871368;
assign addr[13793]= 2004574453;
assign addr[13794]= 2030734582;
assign addr[13795]= 2054318569;
assign addr[13796]= 2075296495;
assign addr[13797]= 2093641749;
assign addr[13798]= 2109331059;
assign addr[13799]= 2122344521;
assign addr[13800]= 2132665626;
assign addr[13801]= 2140281282;
assign addr[13802]= 2145181827;
assign addr[13803]= 2147361045;
assign addr[13804]= 2146816171;
assign addr[13805]= 2143547897;
assign addr[13806]= 2137560369;
assign addr[13807]= 2128861181;
assign addr[13808]= 2117461370;
assign addr[13809]= 2103375398;
assign addr[13810]= 2086621133;
assign addr[13811]= 2067219829;
assign addr[13812]= 2045196100;
assign addr[13813]= 2020577882;
assign addr[13814]= 1993396407;
assign addr[13815]= 1963686155;
assign addr[13816]= 1931484818;
assign addr[13817]= 1896833245;
assign addr[13818]= 1859775393;
assign addr[13819]= 1820358275;
assign addr[13820]= 1778631892;
assign addr[13821]= 1734649179;
assign addr[13822]= 1688465931;
assign addr[13823]= 1640140734;
assign addr[13824]= 1589734894;
assign addr[13825]= 1537312353;
assign addr[13826]= 1482939614;
assign addr[13827]= 1426685652;
assign addr[13828]= 1368621831;
assign addr[13829]= 1308821808;
assign addr[13830]= 1247361445;
assign addr[13831]= 1184318708;
assign addr[13832]= 1119773573;
assign addr[13833]= 1053807919;
assign addr[13834]= 986505429;
assign addr[13835]= 917951481;
assign addr[13836]= 848233042;
assign addr[13837]= 777438554;
assign addr[13838]= 705657826;
assign addr[13839]= 632981917;
assign addr[13840]= 559503022;
assign addr[13841]= 485314355;
assign addr[13842]= 410510029;
assign addr[13843]= 335184940;
assign addr[13844]= 259434643;
assign addr[13845]= 183355234;
assign addr[13846]= 107043224;
assign addr[13847]= 30595422;
assign addr[13848]= -45891193;
assign addr[13849]= -122319591;
assign addr[13850]= -198592817;
assign addr[13851]= -274614114;
assign addr[13852]= -350287041;
assign addr[13853]= -425515602;
assign addr[13854]= -500204365;
assign addr[13855]= -574258580;
assign addr[13856]= -647584304;
assign addr[13857]= -720088517;
assign addr[13858]= -791679244;
assign addr[13859]= -862265664;
assign addr[13860]= -931758235;
assign addr[13861]= -1000068799;
assign addr[13862]= -1067110699;
assign addr[13863]= -1132798888;
assign addr[13864]= -1197050035;
assign addr[13865]= -1259782632;
assign addr[13866]= -1320917099;
assign addr[13867]= -1380375881;
assign addr[13868]= -1438083551;
assign addr[13869]= -1493966902;
assign addr[13870]= -1547955041;
assign addr[13871]= -1599979481;
assign addr[13872]= -1649974225;
assign addr[13873]= -1697875851;
assign addr[13874]= -1743623590;
assign addr[13875]= -1787159411;
assign addr[13876]= -1828428082;
assign addr[13877]= -1867377253;
assign addr[13878]= -1903957513;
assign addr[13879]= -1938122457;
assign addr[13880]= -1969828744;
assign addr[13881]= -1999036154;
assign addr[13882]= -2025707632;
assign addr[13883]= -2049809346;
assign addr[13884]= -2071310720;
assign addr[13885]= -2090184478;
assign addr[13886]= -2106406677;
assign addr[13887]= -2119956737;
assign addr[13888]= -2130817471;
assign addr[13889]= -2138975100;
assign addr[13890]= -2144419275;
assign addr[13891]= -2147143090;
assign addr[13892]= -2147143090;
assign addr[13893]= -2144419275;
assign addr[13894]= -2138975100;
assign addr[13895]= -2130817471;
assign addr[13896]= -2119956737;
assign addr[13897]= -2106406677;
assign addr[13898]= -2090184478;
assign addr[13899]= -2071310720;
assign addr[13900]= -2049809346;
assign addr[13901]= -2025707632;
assign addr[13902]= -1999036154;
assign addr[13903]= -1969828744;
assign addr[13904]= -1938122457;
assign addr[13905]= -1903957513;
assign addr[13906]= -1867377253;
assign addr[13907]= -1828428082;
assign addr[13908]= -1787159411;
assign addr[13909]= -1743623590;
assign addr[13910]= -1697875851;
assign addr[13911]= -1649974225;
assign addr[13912]= -1599979481;
assign addr[13913]= -1547955041;
assign addr[13914]= -1493966902;
assign addr[13915]= -1438083551;
assign addr[13916]= -1380375881;
assign addr[13917]= -1320917099;
assign addr[13918]= -1259782632;
assign addr[13919]= -1197050035;
assign addr[13920]= -1132798888;
assign addr[13921]= -1067110699;
assign addr[13922]= -1000068799;
assign addr[13923]= -931758235;
assign addr[13924]= -862265664;
assign addr[13925]= -791679244;
assign addr[13926]= -720088517;
assign addr[13927]= -647584304;
assign addr[13928]= -574258580;
assign addr[13929]= -500204365;
assign addr[13930]= -425515602;
assign addr[13931]= -350287041;
assign addr[13932]= -274614114;
assign addr[13933]= -198592817;
assign addr[13934]= -122319591;
assign addr[13935]= -45891193;
assign addr[13936]= 30595422;
assign addr[13937]= 107043224;
assign addr[13938]= 183355234;
assign addr[13939]= 259434643;
assign addr[13940]= 335184940;
assign addr[13941]= 410510029;
assign addr[13942]= 485314355;
assign addr[13943]= 559503022;
assign addr[13944]= 632981917;
assign addr[13945]= 705657826;
assign addr[13946]= 777438554;
assign addr[13947]= 848233042;
assign addr[13948]= 917951481;
assign addr[13949]= 986505429;
assign addr[13950]= 1053807919;
assign addr[13951]= 1119773573;
assign addr[13952]= 1184318708;
assign addr[13953]= 1247361445;
assign addr[13954]= 1308821808;
assign addr[13955]= 1368621831;
assign addr[13956]= 1426685652;
assign addr[13957]= 1482939614;
assign addr[13958]= 1537312353;
assign addr[13959]= 1589734894;
assign addr[13960]= 1640140734;
assign addr[13961]= 1688465931;
assign addr[13962]= 1734649179;
assign addr[13963]= 1778631892;
assign addr[13964]= 1820358275;
assign addr[13965]= 1859775393;
assign addr[13966]= 1896833245;
assign addr[13967]= 1931484818;
assign addr[13968]= 1963686155;
assign addr[13969]= 1993396407;
assign addr[13970]= 2020577882;
assign addr[13971]= 2045196100;
assign addr[13972]= 2067219829;
assign addr[13973]= 2086621133;
assign addr[13974]= 2103375398;
assign addr[13975]= 2117461370;
assign addr[13976]= 2128861181;
assign addr[13977]= 2137560369;
assign addr[13978]= 2143547897;
assign addr[13979]= 2146816171;
assign addr[13980]= 2147361045;
assign addr[13981]= 2145181827;
assign addr[13982]= 2140281282;
assign addr[13983]= 2132665626;
assign addr[13984]= 2122344521;
assign addr[13985]= 2109331059;
assign addr[13986]= 2093641749;
assign addr[13987]= 2075296495;
assign addr[13988]= 2054318569;
assign addr[13989]= 2030734582;
assign addr[13990]= 2004574453;
assign addr[13991]= 1975871368;
assign addr[13992]= 1944661739;
assign addr[13993]= 1910985158;
assign addr[13994]= 1874884346;
assign addr[13995]= 1836405100;
assign addr[13996]= 1795596234;
assign addr[13997]= 1752509516;
assign addr[13998]= 1707199606;
assign addr[13999]= 1659723983;
assign addr[14000]= 1610142873;
assign addr[14001]= 1558519173;
assign addr[14002]= 1504918373;
assign addr[14003]= 1449408469;
assign addr[14004]= 1392059879;
assign addr[14005]= 1332945355;
assign addr[14006]= 1272139887;
assign addr[14007]= 1209720613;
assign addr[14008]= 1145766716;
assign addr[14009]= 1080359326;
assign addr[14010]= 1013581418;
assign addr[14011]= 945517704;
assign addr[14012]= 876254528;
assign addr[14013]= 805879757;
assign addr[14014]= 734482665;
assign addr[14015]= 662153826;
assign addr[14016]= 588984994;
assign addr[14017]= 515068990;
assign addr[14018]= 440499581;
assign addr[14019]= 365371365;
assign addr[14020]= 289779648;
assign addr[14021]= 213820322;
assign addr[14022]= 137589750;
assign addr[14023]= 61184634;
assign addr[14024]= -15298099;
assign addr[14025]= -91761426;
assign addr[14026]= -168108346;
assign addr[14027]= -244242007;
assign addr[14028]= -320065829;
assign addr[14029]= -395483624;
assign addr[14030]= -470399716;
assign addr[14031]= -544719071;
assign addr[14032]= -618347408;
assign addr[14033]= -691191324;
assign addr[14034]= -763158411;
assign addr[14035]= -834157373;
assign addr[14036]= -904098143;
assign addr[14037]= -972891995;
assign addr[14038]= -1040451659;
assign addr[14039]= -1106691431;
assign addr[14040]= -1171527280;
assign addr[14041]= -1234876957;
assign addr[14042]= -1296660098;
assign addr[14043]= -1356798326;
assign addr[14044]= -1415215352;
assign addr[14045]= -1471837070;
assign addr[14046]= -1526591649;
assign addr[14047]= -1579409630;
assign addr[14048]= -1630224009;
assign addr[14049]= -1678970324;
assign addr[14050]= -1725586737;
assign addr[14051]= -1770014111;
assign addr[14052]= -1812196087;
assign addr[14053]= -1852079154;
assign addr[14054]= -1889612716;
assign addr[14055]= -1924749160;
assign addr[14056]= -1957443913;
assign addr[14057]= -1987655498;
assign addr[14058]= -2015345591;
assign addr[14059]= -2040479063;
assign addr[14060]= -2063024031;
assign addr[14061]= -2082951896;
assign addr[14062]= -2100237377;
assign addr[14063]= -2114858546;
assign addr[14064]= -2126796855;
assign addr[14065]= -2136037160;
assign addr[14066]= -2142567738;
assign addr[14067]= -2146380306;
assign addr[14068]= -2147470025;
assign addr[14069]= -2145835515;
assign addr[14070]= -2141478848;
assign addr[14071]= -2134405552;
assign addr[14072]= -2124624598;
assign addr[14073]= -2112148396;
assign addr[14074]= -2096992772;
assign addr[14075]= -2079176953;
assign addr[14076]= -2058723538;
assign addr[14077]= -2035658475;
assign addr[14078]= -2010011024;
assign addr[14079]= -1981813720;
assign addr[14080]= -1951102334;
assign addr[14081]= -1917915825;
assign addr[14082]= -1882296293;
assign addr[14083]= -1844288924;
assign addr[14084]= -1803941934;
assign addr[14085]= -1761306505;
assign addr[14086]= -1716436725;
assign addr[14087]= -1669389513;
assign addr[14088]= -1620224553;
assign addr[14089]= -1569004214;
assign addr[14090]= -1515793473;
assign addr[14091]= -1460659832;
assign addr[14092]= -1403673233;
assign addr[14093]= -1344905966;
assign addr[14094]= -1284432584;
assign addr[14095]= -1222329801;
assign addr[14096]= -1158676398;
assign addr[14097]= -1093553126;
assign addr[14098]= -1027042599;
assign addr[14099]= -959229189;
assign addr[14100]= -890198924;
assign addr[14101]= -820039373;
assign addr[14102]= -748839539;
assign addr[14103]= -676689746;
assign addr[14104]= -603681519;
assign addr[14105]= -529907477;
assign addr[14106]= -455461206;
assign addr[14107]= -380437148;
assign addr[14108]= -304930476;
assign addr[14109]= -229036977;
assign addr[14110]= -152852926;
assign addr[14111]= -76474970;
assign addr[14112]= 0;
assign addr[14113]= 76474970;
assign addr[14114]= 152852926;
assign addr[14115]= 229036977;
assign addr[14116]= 304930476;
assign addr[14117]= 380437148;
assign addr[14118]= 455461206;
assign addr[14119]= 529907477;
assign addr[14120]= 603681519;
assign addr[14121]= 676689746;
assign addr[14122]= 748839539;
assign addr[14123]= 820039373;
assign addr[14124]= 890198924;
assign addr[14125]= 959229189;
assign addr[14126]= 1027042599;
assign addr[14127]= 1093553126;
assign addr[14128]= 1158676398;
assign addr[14129]= 1222329801;
assign addr[14130]= 1284432584;
assign addr[14131]= 1344905966;
assign addr[14132]= 1403673233;
assign addr[14133]= 1460659832;
assign addr[14134]= 1515793473;
assign addr[14135]= 1569004214;
assign addr[14136]= 1620224553;
assign addr[14137]= 1669389513;
assign addr[14138]= 1716436725;
assign addr[14139]= 1761306505;
assign addr[14140]= 1803941934;
assign addr[14141]= 1844288924;
assign addr[14142]= 1882296293;
assign addr[14143]= 1917915825;
assign addr[14144]= 1951102334;
assign addr[14145]= 1981813720;
assign addr[14146]= 2010011024;
assign addr[14147]= 2035658475;
assign addr[14148]= 2058723538;
assign addr[14149]= 2079176953;
assign addr[14150]= 2096992772;
assign addr[14151]= 2112148396;
assign addr[14152]= 2124624598;
assign addr[14153]= 2134405552;
assign addr[14154]= 2141478848;
assign addr[14155]= 2145835515;
assign addr[14156]= 2147470025;
assign addr[14157]= 2146380306;
assign addr[14158]= 2142567738;
assign addr[14159]= 2136037160;
assign addr[14160]= 2126796855;
assign addr[14161]= 2114858546;
assign addr[14162]= 2100237377;
assign addr[14163]= 2082951896;
assign addr[14164]= 2063024031;
assign addr[14165]= 2040479063;
assign addr[14166]= 2015345591;
assign addr[14167]= 1987655498;
assign addr[14168]= 1957443913;
assign addr[14169]= 1924749160;
assign addr[14170]= 1889612716;
assign addr[14171]= 1852079154;
assign addr[14172]= 1812196087;
assign addr[14173]= 1770014111;
assign addr[14174]= 1725586737;
assign addr[14175]= 1678970324;
assign addr[14176]= 1630224009;
assign addr[14177]= 1579409630;
assign addr[14178]= 1526591649;
assign addr[14179]= 1471837070;
assign addr[14180]= 1415215352;
assign addr[14181]= 1356798326;
assign addr[14182]= 1296660098;
assign addr[14183]= 1234876957;
assign addr[14184]= 1171527280;
assign addr[14185]= 1106691431;
assign addr[14186]= 1040451659;
assign addr[14187]= 972891995;
assign addr[14188]= 904098143;
assign addr[14189]= 834157373;
assign addr[14190]= 763158411;
assign addr[14191]= 691191324;
assign addr[14192]= 618347408;
assign addr[14193]= 544719071;
assign addr[14194]= 470399716;
assign addr[14195]= 395483624;
assign addr[14196]= 320065829;
assign addr[14197]= 244242007;
assign addr[14198]= 168108346;
assign addr[14199]= 91761426;
assign addr[14200]= 15298099;
assign addr[14201]= -61184634;
assign addr[14202]= -137589750;
assign addr[14203]= -213820322;
assign addr[14204]= -289779648;
assign addr[14205]= -365371365;
assign addr[14206]= -440499581;
assign addr[14207]= -515068990;
assign addr[14208]= -588984994;
assign addr[14209]= -662153826;
assign addr[14210]= -734482665;
assign addr[14211]= -805879757;
assign addr[14212]= -876254528;
assign addr[14213]= -945517704;
assign addr[14214]= -1013581418;
assign addr[14215]= -1080359326;
assign addr[14216]= -1145766716;
assign addr[14217]= -1209720613;
assign addr[14218]= -1272139887;
assign addr[14219]= -1332945355;
assign addr[14220]= -1392059879;
assign addr[14221]= -1449408469;
assign addr[14222]= -1504918373;
assign addr[14223]= -1558519173;
assign addr[14224]= -1610142873;
assign addr[14225]= -1659723983;
assign addr[14226]= -1707199606;
assign addr[14227]= -1752509516;
assign addr[14228]= -1795596234;
assign addr[14229]= -1836405100;
assign addr[14230]= -1874884346;
assign addr[14231]= -1910985158;
assign addr[14232]= -1944661739;
assign addr[14233]= -1975871368;
assign addr[14234]= -2004574453;
assign addr[14235]= -2030734582;
assign addr[14236]= -2054318569;
assign addr[14237]= -2075296495;
assign addr[14238]= -2093641749;
assign addr[14239]= -2109331059;
assign addr[14240]= -2122344521;
assign addr[14241]= -2132665626;
assign addr[14242]= -2140281282;
assign addr[14243]= -2145181827;
assign addr[14244]= -2147361045;
assign addr[14245]= -2146816171;
assign addr[14246]= -2143547897;
assign addr[14247]= -2137560369;
assign addr[14248]= -2128861181;
assign addr[14249]= -2117461370;
assign addr[14250]= -2103375398;
assign addr[14251]= -2086621133;
assign addr[14252]= -2067219829;
assign addr[14253]= -2045196100;
assign addr[14254]= -2020577882;
assign addr[14255]= -1993396407;
assign addr[14256]= -1963686155;
assign addr[14257]= -1931484818;
assign addr[14258]= -1896833245;
assign addr[14259]= -1859775393;
assign addr[14260]= -1820358275;
assign addr[14261]= -1778631892;
assign addr[14262]= -1734649179;
assign addr[14263]= -1688465931;
assign addr[14264]= -1640140734;
assign addr[14265]= -1589734894;
assign addr[14266]= -1537312353;
assign addr[14267]= -1482939614;
assign addr[14268]= -1426685652;
assign addr[14269]= -1368621831;
assign addr[14270]= -1308821808;
assign addr[14271]= -1247361445;
assign addr[14272]= -1184318708;
assign addr[14273]= -1119773573;
assign addr[14274]= -1053807919;
assign addr[14275]= -986505429;
assign addr[14276]= -917951481;
assign addr[14277]= -848233042;
assign addr[14278]= -777438554;
assign addr[14279]= -705657826;
assign addr[14280]= -632981917;
assign addr[14281]= -559503022;
assign addr[14282]= -485314355;
assign addr[14283]= -410510029;
assign addr[14284]= -335184940;
assign addr[14285]= -259434643;
assign addr[14286]= -183355234;
assign addr[14287]= -107043224;
assign addr[14288]= -30595422;
assign addr[14289]= 45891193;
assign addr[14290]= 122319591;
assign addr[14291]= 198592817;
assign addr[14292]= 274614114;
assign addr[14293]= 350287041;
assign addr[14294]= 425515602;
assign addr[14295]= 500204365;
assign addr[14296]= 574258580;
assign addr[14297]= 647584304;
assign addr[14298]= 720088517;
assign addr[14299]= 791679244;
assign addr[14300]= 862265664;
assign addr[14301]= 931758235;
assign addr[14302]= 1000068799;
assign addr[14303]= 1067110699;
assign addr[14304]= 1132798888;
assign addr[14305]= 1197050035;
assign addr[14306]= 1259782632;
assign addr[14307]= 1320917099;
assign addr[14308]= 1380375881;
assign addr[14309]= 1438083551;
assign addr[14310]= 1493966902;
assign addr[14311]= 1547955041;
assign addr[14312]= 1599979481;
assign addr[14313]= 1649974225;
assign addr[14314]= 1697875851;
assign addr[14315]= 1743623590;
assign addr[14316]= 1787159411;
assign addr[14317]= 1828428082;
assign addr[14318]= 1867377253;
assign addr[14319]= 1903957513;
assign addr[14320]= 1938122457;
assign addr[14321]= 1969828744;
assign addr[14322]= 1999036154;
assign addr[14323]= 2025707632;
assign addr[14324]= 2049809346;
assign addr[14325]= 2071310720;
assign addr[14326]= 2090184478;
assign addr[14327]= 2106406677;
assign addr[14328]= 2119956737;
assign addr[14329]= 2130817471;
assign addr[14330]= 2138975100;
assign addr[14331]= 2144419275;
assign addr[14332]= 2147143090;
assign addr[14333]= 2147143090;
assign addr[14334]= 2144419275;
assign addr[14335]= 2138975100;
assign addr[14336]= 2130817471;
assign addr[14337]= 2119956737;
assign addr[14338]= 2106406677;
assign addr[14339]= 2090184478;
assign addr[14340]= 2071310720;
assign addr[14341]= 2049809346;
assign addr[14342]= 2025707632;
assign addr[14343]= 1999036154;
assign addr[14344]= 1969828744;
assign addr[14345]= 1938122457;
assign addr[14346]= 1903957513;
assign addr[14347]= 1867377253;
assign addr[14348]= 1828428082;
assign addr[14349]= 1787159411;
assign addr[14350]= 1743623590;
assign addr[14351]= 1697875851;
assign addr[14352]= 1649974225;
assign addr[14353]= 1599979481;
assign addr[14354]= 1547955041;
assign addr[14355]= 1493966902;
assign addr[14356]= 1438083551;
assign addr[14357]= 1380375881;
assign addr[14358]= 1320917099;
assign addr[14359]= 1259782632;
assign addr[14360]= 1197050035;
assign addr[14361]= 1132798888;
assign addr[14362]= 1067110699;
assign addr[14363]= 1000068799;
assign addr[14364]= 931758235;
assign addr[14365]= 862265664;
assign addr[14366]= 791679244;
assign addr[14367]= 720088517;
assign addr[14368]= 647584304;
assign addr[14369]= 574258580;
assign addr[14370]= 500204365;
assign addr[14371]= 425515602;
assign addr[14372]= 350287041;
assign addr[14373]= 274614114;
assign addr[14374]= 198592817;
assign addr[14375]= 122319591;
assign addr[14376]= 45891193;
assign addr[14377]= -30595422;
assign addr[14378]= -107043224;
assign addr[14379]= -183355234;
assign addr[14380]= -259434643;
assign addr[14381]= -335184940;
assign addr[14382]= -410510029;
assign addr[14383]= -485314355;
assign addr[14384]= -559503022;
assign addr[14385]= -632981917;
assign addr[14386]= -705657826;
assign addr[14387]= -777438554;
assign addr[14388]= -848233042;
assign addr[14389]= -917951481;
assign addr[14390]= -986505429;
assign addr[14391]= -1053807919;
assign addr[14392]= -1119773573;
assign addr[14393]= -1184318708;
assign addr[14394]= -1247361445;
assign addr[14395]= -1308821808;
assign addr[14396]= -1368621831;
assign addr[14397]= -1426685652;
assign addr[14398]= -1482939614;
assign addr[14399]= -1537312353;
assign addr[14400]= -1589734894;
assign addr[14401]= -1640140734;
assign addr[14402]= -1688465931;
assign addr[14403]= -1734649179;
assign addr[14404]= -1778631892;
assign addr[14405]= -1820358275;
assign addr[14406]= -1859775393;
assign addr[14407]= -1896833245;
assign addr[14408]= -1931484818;
assign addr[14409]= -1963686155;
assign addr[14410]= -1993396407;
assign addr[14411]= -2020577882;
assign addr[14412]= -2045196100;
assign addr[14413]= -2067219829;
assign addr[14414]= -2086621133;
assign addr[14415]= -2103375398;
assign addr[14416]= -2117461370;
assign addr[14417]= -2128861181;
assign addr[14418]= -2137560369;
assign addr[14419]= -2143547897;
assign addr[14420]= -2146816171;
assign addr[14421]= -2147361045;
assign addr[14422]= -2145181827;
assign addr[14423]= -2140281282;
assign addr[14424]= -2132665626;
assign addr[14425]= -2122344521;
assign addr[14426]= -2109331059;
assign addr[14427]= -2093641749;
assign addr[14428]= -2075296495;
assign addr[14429]= -2054318569;
assign addr[14430]= -2030734582;
assign addr[14431]= -2004574453;
assign addr[14432]= -1975871368;
assign addr[14433]= -1944661739;
assign addr[14434]= -1910985158;
assign addr[14435]= -1874884346;
assign addr[14436]= -1836405100;
assign addr[14437]= -1795596234;
assign addr[14438]= -1752509516;
assign addr[14439]= -1707199606;
assign addr[14440]= -1659723983;
assign addr[14441]= -1610142873;
assign addr[14442]= -1558519173;
assign addr[14443]= -1504918373;
assign addr[14444]= -1449408469;
assign addr[14445]= -1392059879;
assign addr[14446]= -1332945355;
assign addr[14447]= -1272139887;
assign addr[14448]= -1209720613;
assign addr[14449]= -1145766716;
assign addr[14450]= -1080359326;
assign addr[14451]= -1013581418;
assign addr[14452]= -945517704;
assign addr[14453]= -876254528;
assign addr[14454]= -805879757;
assign addr[14455]= -734482665;
assign addr[14456]= -662153826;
assign addr[14457]= -588984994;
assign addr[14458]= -515068990;
assign addr[14459]= -440499581;
assign addr[14460]= -365371365;
assign addr[14461]= -289779648;
assign addr[14462]= -213820322;
assign addr[14463]= -137589750;
assign addr[14464]= -61184634;
assign addr[14465]= 15298099;
assign addr[14466]= 91761426;
assign addr[14467]= 168108346;
assign addr[14468]= 244242007;
assign addr[14469]= 320065829;
assign addr[14470]= 395483624;
assign addr[14471]= 470399716;
assign addr[14472]= 544719071;
assign addr[14473]= 618347408;
assign addr[14474]= 691191324;
assign addr[14475]= 763158411;
assign addr[14476]= 834157373;
assign addr[14477]= 904098143;
assign addr[14478]= 972891995;
assign addr[14479]= 1040451659;
assign addr[14480]= 1106691431;
assign addr[14481]= 1171527280;
assign addr[14482]= 1234876957;
assign addr[14483]= 1296660098;
assign addr[14484]= 1356798326;
assign addr[14485]= 1415215352;
assign addr[14486]= 1471837070;
assign addr[14487]= 1526591649;
assign addr[14488]= 1579409630;
assign addr[14489]= 1630224009;
assign addr[14490]= 1678970324;
assign addr[14491]= 1725586737;
assign addr[14492]= 1770014111;
assign addr[14493]= 1812196087;
assign addr[14494]= 1852079154;
assign addr[14495]= 1889612716;
assign addr[14496]= 1924749160;
assign addr[14497]= 1957443913;
assign addr[14498]= 1987655498;
assign addr[14499]= 2015345591;
assign addr[14500]= 2040479063;
assign addr[14501]= 2063024031;
assign addr[14502]= 2082951896;
assign addr[14503]= 2100237377;
assign addr[14504]= 2114858546;
assign addr[14505]= 2126796855;
assign addr[14506]= 2136037160;
assign addr[14507]= 2142567738;
assign addr[14508]= 2146380306;
assign addr[14509]= 2147470025;
assign addr[14510]= 2145835515;
assign addr[14511]= 2141478848;
assign addr[14512]= 2134405552;
assign addr[14513]= 2124624598;
assign addr[14514]= 2112148396;
assign addr[14515]= 2096992772;
assign addr[14516]= 2079176953;
assign addr[14517]= 2058723538;
assign addr[14518]= 2035658475;
assign addr[14519]= 2010011024;
assign addr[14520]= 1981813720;
assign addr[14521]= 1951102334;
assign addr[14522]= 1917915825;
assign addr[14523]= 1882296293;
assign addr[14524]= 1844288924;
assign addr[14525]= 1803941934;
assign addr[14526]= 1761306505;
assign addr[14527]= 1716436725;
assign addr[14528]= 1669389513;
assign addr[14529]= 1620224553;
assign addr[14530]= 1569004214;
assign addr[14531]= 1515793473;
assign addr[14532]= 1460659832;
assign addr[14533]= 1403673233;
assign addr[14534]= 1344905966;
assign addr[14535]= 1284432584;
assign addr[14536]= 1222329801;
assign addr[14537]= 1158676398;
assign addr[14538]= 1093553126;
assign addr[14539]= 1027042599;
assign addr[14540]= 959229189;
assign addr[14541]= 890198924;
assign addr[14542]= 820039373;
assign addr[14543]= 748839539;
assign addr[14544]= 676689746;
assign addr[14545]= 603681519;
assign addr[14546]= 529907477;
assign addr[14547]= 455461206;
assign addr[14548]= 380437148;
assign addr[14549]= 304930476;
assign addr[14550]= 229036977;
assign addr[14551]= 152852926;
assign addr[14552]= 76474970;
assign addr[14553]= 0;
assign addr[14554]= -76474970;
assign addr[14555]= -152852926;
assign addr[14556]= -229036977;
assign addr[14557]= -304930476;
assign addr[14558]= -380437148;
assign addr[14559]= -455461206;
assign addr[14560]= -529907477;
assign addr[14561]= -603681519;
assign addr[14562]= -676689746;
assign addr[14563]= -748839539;
assign addr[14564]= -820039373;
assign addr[14565]= -890198924;
assign addr[14566]= -959229189;
assign addr[14567]= -1027042599;
assign addr[14568]= -1093553126;
assign addr[14569]= -1158676398;
assign addr[14570]= -1222329801;
assign addr[14571]= -1284432584;
assign addr[14572]= -1344905966;
assign addr[14573]= -1403673233;
assign addr[14574]= -1460659832;
assign addr[14575]= -1515793473;
assign addr[14576]= -1569004214;
assign addr[14577]= -1620224553;
assign addr[14578]= -1669389513;
assign addr[14579]= -1716436725;
assign addr[14580]= -1761306505;
assign addr[14581]= -1803941934;
assign addr[14582]= -1844288924;
assign addr[14583]= -1882296293;
assign addr[14584]= -1917915825;
assign addr[14585]= -1951102334;
assign addr[14586]= -1981813720;
assign addr[14587]= -2010011024;
assign addr[14588]= -2035658475;
assign addr[14589]= -2058723538;
assign addr[14590]= -2079176953;
assign addr[14591]= -2096992772;
assign addr[14592]= -2112148396;
assign addr[14593]= -2124624598;
assign addr[14594]= -2134405552;
assign addr[14595]= -2141478848;
assign addr[14596]= -2145835515;
assign addr[14597]= -2147470025;
assign addr[14598]= -2146380306;
assign addr[14599]= -2142567738;
assign addr[14600]= -2136037160;
assign addr[14601]= -2126796855;
assign addr[14602]= -2114858546;
assign addr[14603]= -2100237377;
assign addr[14604]= -2082951896;
assign addr[14605]= -2063024031;
assign addr[14606]= -2040479063;
assign addr[14607]= -2015345591;
assign addr[14608]= -1987655498;
assign addr[14609]= -1957443913;
assign addr[14610]= -1924749160;
assign addr[14611]= -1889612716;
assign addr[14612]= -1852079154;
assign addr[14613]= -1812196087;
assign addr[14614]= -1770014111;
assign addr[14615]= -1725586737;
assign addr[14616]= -1678970324;
assign addr[14617]= -1630224009;
assign addr[14618]= -1579409630;
assign addr[14619]= -1526591649;
assign addr[14620]= -1471837070;
assign addr[14621]= -1415215352;
assign addr[14622]= -1356798326;
assign addr[14623]= -1296660098;
assign addr[14624]= -1234876957;
assign addr[14625]= -1171527280;
assign addr[14626]= -1106691431;
assign addr[14627]= -1040451659;
assign addr[14628]= -972891995;
assign addr[14629]= -904098143;
assign addr[14630]= -834157373;
assign addr[14631]= -763158411;
assign addr[14632]= -691191324;
assign addr[14633]= -618347408;
assign addr[14634]= -544719071;
assign addr[14635]= -470399716;
assign addr[14636]= -395483624;
assign addr[14637]= -320065829;
assign addr[14638]= -244242007;
assign addr[14639]= -168108346;
assign addr[14640]= -91761426;
assign addr[14641]= -15298099;
assign addr[14642]= 61184634;
assign addr[14643]= 137589750;
assign addr[14644]= 213820322;
assign addr[14645]= 289779648;
assign addr[14646]= 365371365;
assign addr[14647]= 440499581;
assign addr[14648]= 515068990;
assign addr[14649]= 588984994;
assign addr[14650]= 662153826;
assign addr[14651]= 734482665;
assign addr[14652]= 805879757;
assign addr[14653]= 876254528;
assign addr[14654]= 945517704;
assign addr[14655]= 1013581418;
assign addr[14656]= 1080359326;
assign addr[14657]= 1145766716;
assign addr[14658]= 1209720613;
assign addr[14659]= 1272139887;
assign addr[14660]= 1332945355;
assign addr[14661]= 1392059879;
assign addr[14662]= 1449408469;
assign addr[14663]= 1504918373;
assign addr[14664]= 1558519173;
assign addr[14665]= 1610142873;
assign addr[14666]= 1659723983;
assign addr[14667]= 1707199606;
assign addr[14668]= 1752509516;
assign addr[14669]= 1795596234;
assign addr[14670]= 1836405100;
assign addr[14671]= 1874884346;
assign addr[14672]= 1910985158;
assign addr[14673]= 1944661739;
assign addr[14674]= 1975871368;
assign addr[14675]= 2004574453;
assign addr[14676]= 2030734582;
assign addr[14677]= 2054318569;
assign addr[14678]= 2075296495;
assign addr[14679]= 2093641749;
assign addr[14680]= 2109331059;
assign addr[14681]= 2122344521;
assign addr[14682]= 2132665626;
assign addr[14683]= 2140281282;
assign addr[14684]= 2145181827;
assign addr[14685]= 2147361045;
assign addr[14686]= 2146816171;
assign addr[14687]= 2143547897;
assign addr[14688]= 2137560369;
assign addr[14689]= 2128861181;
assign addr[14690]= 2117461370;
assign addr[14691]= 2103375398;
assign addr[14692]= 2086621133;
assign addr[14693]= 2067219829;
assign addr[14694]= 2045196100;
assign addr[14695]= 2020577882;
assign addr[14696]= 1993396407;
assign addr[14697]= 1963686155;
assign addr[14698]= 1931484818;
assign addr[14699]= 1896833245;
assign addr[14700]= 1859775393;
assign addr[14701]= 1820358275;
assign addr[14702]= 1778631892;
assign addr[14703]= 1734649179;
assign addr[14704]= 1688465931;
assign addr[14705]= 1640140734;
assign addr[14706]= 1589734894;
assign addr[14707]= 1537312353;
assign addr[14708]= 1482939614;
assign addr[14709]= 1426685652;
assign addr[14710]= 1368621831;
assign addr[14711]= 1308821808;
assign addr[14712]= 1247361445;
assign addr[14713]= 1184318708;
assign addr[14714]= 1119773573;
assign addr[14715]= 1053807919;
assign addr[14716]= 986505429;
assign addr[14717]= 917951481;
assign addr[14718]= 848233042;
assign addr[14719]= 777438554;
assign addr[14720]= 705657826;
assign addr[14721]= 632981917;
assign addr[14722]= 559503022;
assign addr[14723]= 485314355;
assign addr[14724]= 410510029;
assign addr[14725]= 335184940;
assign addr[14726]= 259434643;
assign addr[14727]= 183355234;
assign addr[14728]= 107043224;
assign addr[14729]= 30595422;
assign addr[14730]= -45891193;
assign addr[14731]= -122319591;
assign addr[14732]= -198592817;
assign addr[14733]= -274614114;
assign addr[14734]= -350287041;
assign addr[14735]= -425515602;
assign addr[14736]= -500204365;
assign addr[14737]= -574258580;
assign addr[14738]= -647584304;
assign addr[14739]= -720088517;
assign addr[14740]= -791679244;
assign addr[14741]= -862265664;
assign addr[14742]= -931758235;
assign addr[14743]= -1000068799;
assign addr[14744]= -1067110699;
assign addr[14745]= -1132798888;
assign addr[14746]= -1197050035;
assign addr[14747]= -1259782632;
assign addr[14748]= -1320917099;
assign addr[14749]= -1380375881;
assign addr[14750]= -1438083551;
assign addr[14751]= -1493966902;
assign addr[14752]= -1547955041;
assign addr[14753]= -1599979481;
assign addr[14754]= -1649974225;
assign addr[14755]= -1697875851;
assign addr[14756]= -1743623590;
assign addr[14757]= -1787159411;
assign addr[14758]= -1828428082;
assign addr[14759]= -1867377253;
assign addr[14760]= -1903957513;
assign addr[14761]= -1938122457;
assign addr[14762]= -1969828744;
assign addr[14763]= -1999036154;
assign addr[14764]= -2025707632;
assign addr[14765]= -2049809346;
assign addr[14766]= -2071310720;
assign addr[14767]= -2090184478;
assign addr[14768]= -2106406677;
assign addr[14769]= -2119956737;
assign addr[14770]= -2130817471;
assign addr[14771]= -2138975100;
assign addr[14772]= -2144419275;
assign addr[14773]= -2147143090;
assign addr[14774]= -2147143090;
assign addr[14775]= -2144419275;
assign addr[14776]= -2138975100;
assign addr[14777]= -2130817471;
assign addr[14778]= -2119956737;
assign addr[14779]= -2106406677;
assign addr[14780]= -2090184478;
assign addr[14781]= -2071310720;
assign addr[14782]= -2049809346;
assign addr[14783]= -2025707632;
assign addr[14784]= -1999036154;
assign addr[14785]= -1969828744;
assign addr[14786]= -1938122457;
assign addr[14787]= -1903957513;
assign addr[14788]= -1867377253;
assign addr[14789]= -1828428082;
assign addr[14790]= -1787159411;
assign addr[14791]= -1743623590;
assign addr[14792]= -1697875851;
assign addr[14793]= -1649974225;
assign addr[14794]= -1599979481;
assign addr[14795]= -1547955041;
assign addr[14796]= -1493966902;
assign addr[14797]= -1438083551;
assign addr[14798]= -1380375881;
assign addr[14799]= -1320917099;
assign addr[14800]= -1259782632;
assign addr[14801]= -1197050035;
assign addr[14802]= -1132798888;
assign addr[14803]= -1067110699;
assign addr[14804]= -1000068799;
assign addr[14805]= -931758235;
assign addr[14806]= -862265664;
assign addr[14807]= -791679244;
assign addr[14808]= -720088517;
assign addr[14809]= -647584304;
assign addr[14810]= -574258580;
assign addr[14811]= -500204365;
assign addr[14812]= -425515602;
assign addr[14813]= -350287041;
assign addr[14814]= -274614114;
assign addr[14815]= -198592817;
assign addr[14816]= -122319591;
assign addr[14817]= -45891193;
assign addr[14818]= 30595422;
assign addr[14819]= 107043224;
assign addr[14820]= 183355234;
assign addr[14821]= 259434643;
assign addr[14822]= 335184940;
assign addr[14823]= 410510029;
assign addr[14824]= 485314355;
assign addr[14825]= 559503022;
assign addr[14826]= 632981917;
assign addr[14827]= 705657826;
assign addr[14828]= 777438554;
assign addr[14829]= 848233042;
assign addr[14830]= 917951481;
assign addr[14831]= 986505429;
assign addr[14832]= 1053807919;
assign addr[14833]= 1119773573;
assign addr[14834]= 1184318708;
assign addr[14835]= 1247361445;
assign addr[14836]= 1308821808;
assign addr[14837]= 1368621831;
assign addr[14838]= 1426685652;
assign addr[14839]= 1482939614;
assign addr[14840]= 1537312353;
assign addr[14841]= 1589734894;
assign addr[14842]= 1640140734;
assign addr[14843]= 1688465931;
assign addr[14844]= 1734649179;
assign addr[14845]= 1778631892;
assign addr[14846]= 1820358275;
assign addr[14847]= 1859775393;
assign addr[14848]= 1896833245;
assign addr[14849]= 1931484818;
assign addr[14850]= 1963686155;
assign addr[14851]= 1993396407;
assign addr[14852]= 2020577882;
assign addr[14853]= 2045196100;
assign addr[14854]= 2067219829;
assign addr[14855]= 2086621133;
assign addr[14856]= 2103375398;
assign addr[14857]= 2117461370;
assign addr[14858]= 2128861181;
assign addr[14859]= 2137560369;
assign addr[14860]= 2143547897;
assign addr[14861]= 2146816171;
assign addr[14862]= 2147361045;
assign addr[14863]= 2145181827;
assign addr[14864]= 2140281282;
assign addr[14865]= 2132665626;
assign addr[14866]= 2122344521;
assign addr[14867]= 2109331059;
assign addr[14868]= 2093641749;
assign addr[14869]= 2075296495;
assign addr[14870]= 2054318569;
assign addr[14871]= 2030734582;
assign addr[14872]= 2004574453;
assign addr[14873]= 1975871368;
assign addr[14874]= 1944661739;
assign addr[14875]= 1910985158;
assign addr[14876]= 1874884346;
assign addr[14877]= 1836405100;
assign addr[14878]= 1795596234;
assign addr[14879]= 1752509516;
assign addr[14880]= 1707199606;
assign addr[14881]= 1659723983;
assign addr[14882]= 1610142873;
assign addr[14883]= 1558519173;
assign addr[14884]= 1504918373;
assign addr[14885]= 1449408469;
assign addr[14886]= 1392059879;
assign addr[14887]= 1332945355;
assign addr[14888]= 1272139887;
assign addr[14889]= 1209720613;
assign addr[14890]= 1145766716;
assign addr[14891]= 1080359326;
assign addr[14892]= 1013581418;
assign addr[14893]= 945517704;
assign addr[14894]= 876254528;
assign addr[14895]= 805879757;
assign addr[14896]= 734482665;
assign addr[14897]= 662153826;
assign addr[14898]= 588984994;
assign addr[14899]= 515068990;
assign addr[14900]= 440499581;
assign addr[14901]= 365371365;
assign addr[14902]= 289779648;
assign addr[14903]= 213820322;
assign addr[14904]= 137589750;
assign addr[14905]= 61184634;
assign addr[14906]= -15298099;
assign addr[14907]= -91761426;
assign addr[14908]= -168108346;
assign addr[14909]= -244242007;
assign addr[14910]= -320065829;
assign addr[14911]= -395483624;
assign addr[14912]= -470399716;
assign addr[14913]= -544719071;
assign addr[14914]= -618347408;
assign addr[14915]= -691191324;
assign addr[14916]= -763158411;
assign addr[14917]= -834157373;
assign addr[14918]= -904098143;
assign addr[14919]= -972891995;
assign addr[14920]= -1040451659;
assign addr[14921]= -1106691431;
assign addr[14922]= -1171527280;
assign addr[14923]= -1234876957;
assign addr[14924]= -1296660098;
assign addr[14925]= -1356798326;
assign addr[14926]= -1415215352;
assign addr[14927]= -1471837070;
assign addr[14928]= -1526591649;
assign addr[14929]= -1579409630;
assign addr[14930]= -1630224009;
assign addr[14931]= -1678970324;
assign addr[14932]= -1725586737;
assign addr[14933]= -1770014111;
assign addr[14934]= -1812196087;
assign addr[14935]= -1852079154;
assign addr[14936]= -1889612716;
assign addr[14937]= -1924749160;
assign addr[14938]= -1957443913;
assign addr[14939]= -1987655498;
assign addr[14940]= -2015345591;
assign addr[14941]= -2040479063;
assign addr[14942]= -2063024031;
assign addr[14943]= -2082951896;
assign addr[14944]= -2100237377;
assign addr[14945]= -2114858546;
assign addr[14946]= -2126796855;
assign addr[14947]= -2136037160;
assign addr[14948]= -2142567738;
assign addr[14949]= -2146380306;
assign addr[14950]= -2147470025;
assign addr[14951]= -2145835515;
assign addr[14952]= -2141478848;
assign addr[14953]= -2134405552;
assign addr[14954]= -2124624598;
assign addr[14955]= -2112148396;
assign addr[14956]= -2096992772;
assign addr[14957]= -2079176953;
assign addr[14958]= -2058723538;
assign addr[14959]= -2035658475;
assign addr[14960]= -2010011024;
assign addr[14961]= -1981813720;
assign addr[14962]= -1951102334;
assign addr[14963]= -1917915825;
assign addr[14964]= -1882296293;
assign addr[14965]= -1844288924;
assign addr[14966]= -1803941934;
assign addr[14967]= -1761306505;
assign addr[14968]= -1716436725;
assign addr[14969]= -1669389513;
assign addr[14970]= -1620224553;
assign addr[14971]= -1569004214;
assign addr[14972]= -1515793473;
assign addr[14973]= -1460659832;
assign addr[14974]= -1403673233;
assign addr[14975]= -1344905966;
assign addr[14976]= -1284432584;
assign addr[14977]= -1222329801;
assign addr[14978]= -1158676398;
assign addr[14979]= -1093553126;
assign addr[14980]= -1027042599;
assign addr[14981]= -959229189;
assign addr[14982]= -890198924;
assign addr[14983]= -820039373;
assign addr[14984]= -748839539;
assign addr[14985]= -676689746;
assign addr[14986]= -603681519;
assign addr[14987]= -529907477;
assign addr[14988]= -455461206;
assign addr[14989]= -380437148;
assign addr[14990]= -304930476;
assign addr[14991]= -229036977;
assign addr[14992]= -152852926;
assign addr[14993]= -76474970;
assign addr[14994]= 0;
assign addr[14995]= 76474970;
assign addr[14996]= 152852926;
assign addr[14997]= 229036977;
assign addr[14998]= 304930476;
assign addr[14999]= 380437148;
assign addr[15000]= 455461206;
assign addr[15001]= 529907477;
assign addr[15002]= 603681519;
assign addr[15003]= 676689746;
assign addr[15004]= 748839539;
assign addr[15005]= 820039373;
assign addr[15006]= 890198924;
assign addr[15007]= 959229189;
assign addr[15008]= 1027042599;
assign addr[15009]= 1093553126;
assign addr[15010]= 1158676398;
assign addr[15011]= 1222329801;
assign addr[15012]= 1284432584;
assign addr[15013]= 1344905966;
assign addr[15014]= 1403673233;
assign addr[15015]= 1460659832;
assign addr[15016]= 1515793473;
assign addr[15017]= 1569004214;
assign addr[15018]= 1620224553;
assign addr[15019]= 1669389513;
assign addr[15020]= 1716436725;
assign addr[15021]= 1761306505;
assign addr[15022]= 1803941934;
assign addr[15023]= 1844288924;
assign addr[15024]= 1882296293;
assign addr[15025]= 1917915825;
assign addr[15026]= 1951102334;
assign addr[15027]= 1981813720;
assign addr[15028]= 2010011024;
assign addr[15029]= 2035658475;
assign addr[15030]= 2058723538;
assign addr[15031]= 2079176953;
assign addr[15032]= 2096992772;
assign addr[15033]= 2112148396;
assign addr[15034]= 2124624598;
assign addr[15035]= 2134405552;
assign addr[15036]= 2141478848;
assign addr[15037]= 2145835515;
assign addr[15038]= 2147470025;
assign addr[15039]= 2146380306;
assign addr[15040]= 2142567738;
assign addr[15041]= 2136037160;
assign addr[15042]= 2126796855;
assign addr[15043]= 2114858546;
assign addr[15044]= 2100237377;
assign addr[15045]= 2082951896;
assign addr[15046]= 2063024031;
assign addr[15047]= 2040479063;
assign addr[15048]= 2015345591;
assign addr[15049]= 1987655498;
assign addr[15050]= 1957443913;
assign addr[15051]= 1924749160;
assign addr[15052]= 1889612716;
assign addr[15053]= 1852079154;
assign addr[15054]= 1812196087;
assign addr[15055]= 1770014111;
assign addr[15056]= 1725586737;
assign addr[15057]= 1678970324;
assign addr[15058]= 1630224009;
assign addr[15059]= 1579409630;
assign addr[15060]= 1526591649;
assign addr[15061]= 1471837070;
assign addr[15062]= 1415215352;
assign addr[15063]= 1356798326;
assign addr[15064]= 1296660098;
assign addr[15065]= 1234876957;
assign addr[15066]= 1171527280;
assign addr[15067]= 1106691431;
assign addr[15068]= 1040451659;
assign addr[15069]= 972891995;
assign addr[15070]= 904098143;
assign addr[15071]= 834157373;
assign addr[15072]= 763158411;
assign addr[15073]= 691191324;
assign addr[15074]= 618347408;
assign addr[15075]= 544719071;
assign addr[15076]= 470399716;
assign addr[15077]= 395483624;
assign addr[15078]= 320065829;
assign addr[15079]= 244242007;
assign addr[15080]= 168108346;
assign addr[15081]= 91761426;
assign addr[15082]= 15298099;
assign addr[15083]= -61184634;
assign addr[15084]= -137589750;
assign addr[15085]= -213820322;
assign addr[15086]= -289779648;
assign addr[15087]= -365371365;
assign addr[15088]= -440499581;
assign addr[15089]= -515068990;
assign addr[15090]= -588984994;
assign addr[15091]= -662153826;
assign addr[15092]= -734482665;
assign addr[15093]= -805879757;
assign addr[15094]= -876254528;
assign addr[15095]= -945517704;
assign addr[15096]= -1013581418;
assign addr[15097]= -1080359326;
assign addr[15098]= -1145766716;
assign addr[15099]= -1209720613;
assign addr[15100]= -1272139887;
assign addr[15101]= -1332945355;
assign addr[15102]= -1392059879;
assign addr[15103]= -1449408469;
assign addr[15104]= -1504918373;
assign addr[15105]= -1558519173;
assign addr[15106]= -1610142873;
assign addr[15107]= -1659723983;
assign addr[15108]= -1707199606;
assign addr[15109]= -1752509516;
assign addr[15110]= -1795596234;
assign addr[15111]= -1836405100;
assign addr[15112]= -1874884346;
assign addr[15113]= -1910985158;
assign addr[15114]= -1944661739;
assign addr[15115]= -1975871368;
assign addr[15116]= -2004574453;
assign addr[15117]= -2030734582;
assign addr[15118]= -2054318569;
assign addr[15119]= -2075296495;
assign addr[15120]= -2093641749;
assign addr[15121]= -2109331059;
assign addr[15122]= -2122344521;
assign addr[15123]= -2132665626;
assign addr[15124]= -2140281282;
assign addr[15125]= -2145181827;
assign addr[15126]= -2147361045;
assign addr[15127]= -2146816171;
assign addr[15128]= -2143547897;
assign addr[15129]= -2137560369;
assign addr[15130]= -2128861181;
assign addr[15131]= -2117461370;
assign addr[15132]= -2103375398;
assign addr[15133]= -2086621133;
assign addr[15134]= -2067219829;
assign addr[15135]= -2045196100;
assign addr[15136]= -2020577882;
assign addr[15137]= -1993396407;
assign addr[15138]= -1963686155;
assign addr[15139]= -1931484818;
assign addr[15140]= -1896833245;
assign addr[15141]= -1859775393;
assign addr[15142]= -1820358275;
assign addr[15143]= -1778631892;
assign addr[15144]= -1734649179;
assign addr[15145]= -1688465931;
assign addr[15146]= -1640140734;
assign addr[15147]= -1589734894;
assign addr[15148]= -1537312353;
assign addr[15149]= -1482939614;
assign addr[15150]= -1426685652;
assign addr[15151]= -1368621831;
assign addr[15152]= -1308821808;
assign addr[15153]= -1247361445;
assign addr[15154]= -1184318708;
assign addr[15155]= -1119773573;
assign addr[15156]= -1053807919;
assign addr[15157]= -986505429;
assign addr[15158]= -917951481;
assign addr[15159]= -848233042;
assign addr[15160]= -777438554;
assign addr[15161]= -705657826;
assign addr[15162]= -632981917;
assign addr[15163]= -559503022;
assign addr[15164]= -485314355;
assign addr[15165]= -410510029;
assign addr[15166]= -335184940;
assign addr[15167]= -259434643;
assign addr[15168]= -183355234;
assign addr[15169]= -107043224;
assign addr[15170]= -30595422;
assign addr[15171]= 45891193;
assign addr[15172]= 122319591;
assign addr[15173]= 198592817;
assign addr[15174]= 274614114;
assign addr[15175]= 350287041;
assign addr[15176]= 425515602;
assign addr[15177]= 500204365;
assign addr[15178]= 574258580;
assign addr[15179]= 647584304;
assign addr[15180]= 720088517;
assign addr[15181]= 791679244;
assign addr[15182]= 862265664;
assign addr[15183]= 931758235;
assign addr[15184]= 1000068799;
assign addr[15185]= 1067110699;
assign addr[15186]= 1132798888;
assign addr[15187]= 1197050035;
assign addr[15188]= 1259782632;
assign addr[15189]= 1320917099;
assign addr[15190]= 1380375881;
assign addr[15191]= 1438083551;
assign addr[15192]= 1493966902;
assign addr[15193]= 1547955041;
assign addr[15194]= 1599979481;
assign addr[15195]= 1649974225;
assign addr[15196]= 1697875851;
assign addr[15197]= 1743623590;
assign addr[15198]= 1787159411;
assign addr[15199]= 1828428082;
assign addr[15200]= 1867377253;
assign addr[15201]= 1903957513;
assign addr[15202]= 1938122457;
assign addr[15203]= 1969828744;
assign addr[15204]= 1999036154;
assign addr[15205]= 2025707632;
assign addr[15206]= 2049809346;
assign addr[15207]= 2071310720;
assign addr[15208]= 2090184478;
assign addr[15209]= 2106406677;
assign addr[15210]= 2119956737;
assign addr[15211]= 2130817471;
assign addr[15212]= 2138975100;
assign addr[15213]= 2144419275;
assign addr[15214]= 2147143090;
assign addr[15215]= 2147143090;
assign addr[15216]= 2144419275;
assign addr[15217]= 2138975100;
assign addr[15218]= 2130817471;
assign addr[15219]= 2119956737;
assign addr[15220]= 2106406677;
assign addr[15221]= 2090184478;
assign addr[15222]= 2071310720;
assign addr[15223]= 2049809346;
assign addr[15224]= 2025707632;
assign addr[15225]= 1999036154;
assign addr[15226]= 1969828744;
assign addr[15227]= 1938122457;
assign addr[15228]= 1903957513;
assign addr[15229]= 1867377253;
assign addr[15230]= 1828428082;
assign addr[15231]= 1787159411;
assign addr[15232]= 1743623590;
assign addr[15233]= 1697875851;
assign addr[15234]= 1649974225;
assign addr[15235]= 1599979481;
assign addr[15236]= 1547955041;
assign addr[15237]= 1493966902;
assign addr[15238]= 1438083551;
assign addr[15239]= 1380375881;
assign addr[15240]= 1320917099;
assign addr[15241]= 1259782632;
assign addr[15242]= 1197050035;
assign addr[15243]= 1132798888;
assign addr[15244]= 1067110699;
assign addr[15245]= 1000068799;
assign addr[15246]= 931758235;
assign addr[15247]= 862265664;
assign addr[15248]= 791679244;
assign addr[15249]= 720088517;
assign addr[15250]= 647584304;
assign addr[15251]= 574258580;
assign addr[15252]= 500204365;
assign addr[15253]= 425515602;
assign addr[15254]= 350287041;
assign addr[15255]= 274614114;
assign addr[15256]= 198592817;
assign addr[15257]= 122319591;
assign addr[15258]= 45891193;
assign addr[15259]= -30595422;
assign addr[15260]= -107043224;
assign addr[15261]= -183355234;
assign addr[15262]= -259434643;
assign addr[15263]= -335184940;
assign addr[15264]= -410510029;
assign addr[15265]= -485314355;
assign addr[15266]= -559503022;
assign addr[15267]= -632981917;
assign addr[15268]= -705657826;
assign addr[15269]= -777438554;
assign addr[15270]= -848233042;
assign addr[15271]= -917951481;
assign addr[15272]= -986505429;
assign addr[15273]= -1053807919;
assign addr[15274]= -1119773573;
assign addr[15275]= -1184318708;
assign addr[15276]= -1247361445;
assign addr[15277]= -1308821808;
assign addr[15278]= -1368621831;
assign addr[15279]= -1426685652;
assign addr[15280]= -1482939614;
assign addr[15281]= -1537312353;
assign addr[15282]= -1589734894;
assign addr[15283]= -1640140734;
assign addr[15284]= -1688465931;
assign addr[15285]= -1734649179;
assign addr[15286]= -1778631892;
assign addr[15287]= -1820358275;
assign addr[15288]= -1859775393;
assign addr[15289]= -1896833245;
assign addr[15290]= -1931484818;
assign addr[15291]= -1963686155;
assign addr[15292]= -1993396407;
assign addr[15293]= -2020577882;
assign addr[15294]= -2045196100;
assign addr[15295]= -2067219829;
assign addr[15296]= -2086621133;
assign addr[15297]= -2103375398;
assign addr[15298]= -2117461370;
assign addr[15299]= -2128861181;
assign addr[15300]= -2137560369;
assign addr[15301]= -2143547897;
assign addr[15302]= -2146816171;
assign addr[15303]= -2147361045;
assign addr[15304]= -2145181827;
assign addr[15305]= -2140281282;
assign addr[15306]= -2132665626;
assign addr[15307]= -2122344521;
assign addr[15308]= -2109331059;
assign addr[15309]= -2093641749;
assign addr[15310]= -2075296495;
assign addr[15311]= -2054318569;
assign addr[15312]= -2030734582;
assign addr[15313]= -2004574453;
assign addr[15314]= -1975871368;
assign addr[15315]= -1944661739;
assign addr[15316]= -1910985158;
assign addr[15317]= -1874884346;
assign addr[15318]= -1836405100;
assign addr[15319]= -1795596234;
assign addr[15320]= -1752509516;
assign addr[15321]= -1707199606;
assign addr[15322]= -1659723983;
assign addr[15323]= -1610142873;
assign addr[15324]= -1558519173;
assign addr[15325]= -1504918373;
assign addr[15326]= -1449408469;
assign addr[15327]= -1392059879;
assign addr[15328]= -1332945355;
assign addr[15329]= -1272139887;
assign addr[15330]= -1209720613;
assign addr[15331]= -1145766716;
assign addr[15332]= -1080359326;
assign addr[15333]= -1013581418;
assign addr[15334]= -945517704;
assign addr[15335]= -876254528;
assign addr[15336]= -805879757;
assign addr[15337]= -734482665;
assign addr[15338]= -662153826;
assign addr[15339]= -588984994;
assign addr[15340]= -515068990;
assign addr[15341]= -440499581;
assign addr[15342]= -365371365;
assign addr[15343]= -289779648;
assign addr[15344]= -213820322;
assign addr[15345]= -137589750;
assign addr[15346]= -61184634;
assign addr[15347]= 15298099;
assign addr[15348]= 91761426;
assign addr[15349]= 168108346;
assign addr[15350]= 244242007;
assign addr[15351]= 320065829;
assign addr[15352]= 395483624;
assign addr[15353]= 470399716;
assign addr[15354]= 544719071;
assign addr[15355]= 618347408;
assign addr[15356]= 691191324;
assign addr[15357]= 763158411;
assign addr[15358]= 834157373;
assign addr[15359]= 904098143;
assign addr[15360]= 972891995;
assign addr[15361]= 1040451659;
assign addr[15362]= 1106691431;
assign addr[15363]= 1171527280;
assign addr[15364]= 1234876957;
assign addr[15365]= 1296660098;
assign addr[15366]= 1356798326;
assign addr[15367]= 1415215352;
assign addr[15368]= 1471837070;
assign addr[15369]= 1526591649;
assign addr[15370]= 1579409630;
assign addr[15371]= 1630224009;
assign addr[15372]= 1678970324;
assign addr[15373]= 1725586737;
assign addr[15374]= 1770014111;
assign addr[15375]= 1812196087;
assign addr[15376]= 1852079154;
assign addr[15377]= 1889612716;
assign addr[15378]= 1924749160;
assign addr[15379]= 1957443913;
assign addr[15380]= 1987655498;
assign addr[15381]= 2015345591;
assign addr[15382]= 2040479063;
assign addr[15383]= 2063024031;
assign addr[15384]= 2082951896;
assign addr[15385]= 2100237377;
assign addr[15386]= 2114858546;
assign addr[15387]= 2126796855;
assign addr[15388]= 2136037160;
assign addr[15389]= 2142567738;
assign addr[15390]= 2146380306;
assign addr[15391]= 2147470025;
assign addr[15392]= 2145835515;
assign addr[15393]= 2141478848;
assign addr[15394]= 2134405552;
assign addr[15395]= 2124624598;
assign addr[15396]= 2112148396;
assign addr[15397]= 2096992772;
assign addr[15398]= 2079176953;
assign addr[15399]= 2058723538;
assign addr[15400]= 2035658475;
assign addr[15401]= 2010011024;
assign addr[15402]= 1981813720;
assign addr[15403]= 1951102334;
assign addr[15404]= 1917915825;
assign addr[15405]= 1882296293;
assign addr[15406]= 1844288924;
assign addr[15407]= 1803941934;
assign addr[15408]= 1761306505;
assign addr[15409]= 1716436725;
assign addr[15410]= 1669389513;
assign addr[15411]= 1620224553;
assign addr[15412]= 1569004214;
assign addr[15413]= 1515793473;
assign addr[15414]= 1460659832;
assign addr[15415]= 1403673233;
assign addr[15416]= 1344905966;
assign addr[15417]= 1284432584;
assign addr[15418]= 1222329801;
assign addr[15419]= 1158676398;
assign addr[15420]= 1093553126;
assign addr[15421]= 1027042599;
assign addr[15422]= 959229189;
assign addr[15423]= 890198924;
assign addr[15424]= 820039373;
assign addr[15425]= 748839539;
assign addr[15426]= 676689746;
assign addr[15427]= 603681519;
assign addr[15428]= 529907477;
assign addr[15429]= 455461206;
assign addr[15430]= 380437148;
assign addr[15431]= 304930476;
assign addr[15432]= 229036977;
assign addr[15433]= 152852926;
assign addr[15434]= 76474970;
assign addr[15435]= 0;
assign addr[15436]= -76474970;
assign addr[15437]= -152852926;
assign addr[15438]= -229036977;
assign addr[15439]= -304930476;
assign addr[15440]= -380437148;
assign addr[15441]= -455461206;
assign addr[15442]= -529907477;
assign addr[15443]= -603681519;
assign addr[15444]= -676689746;
assign addr[15445]= -748839539;
assign addr[15446]= -820039373;
assign addr[15447]= -890198924;
assign addr[15448]= -959229189;
assign addr[15449]= -1027042599;
assign addr[15450]= -1093553126;
assign addr[15451]= -1158676398;
assign addr[15452]= -1222329801;
assign addr[15453]= -1284432584;
assign addr[15454]= -1344905966;
assign addr[15455]= -1403673233;
assign addr[15456]= -1460659832;
assign addr[15457]= -1515793473;
assign addr[15458]= -1569004214;
assign addr[15459]= -1620224553;
assign addr[15460]= -1669389513;
assign addr[15461]= -1716436725;
assign addr[15462]= -1761306505;
assign addr[15463]= -1803941934;
assign addr[15464]= -1844288924;
assign addr[15465]= -1882296293;
assign addr[15466]= -1917915825;
assign addr[15467]= -1951102334;
assign addr[15468]= -1981813720;
assign addr[15469]= -2010011024;
assign addr[15470]= -2035658475;
assign addr[15471]= -2058723538;
assign addr[15472]= -2079176953;
assign addr[15473]= -2096992772;
assign addr[15474]= -2112148396;
assign addr[15475]= -2124624598;
assign addr[15476]= -2134405552;
assign addr[15477]= -2141478848;
assign addr[15478]= -2145835515;
assign addr[15479]= -2147470025;
assign addr[15480]= -2146380306;
assign addr[15481]= -2142567738;
assign addr[15482]= -2136037160;
assign addr[15483]= -2126796855;
assign addr[15484]= -2114858546;
assign addr[15485]= -2100237377;
assign addr[15486]= -2082951896;
assign addr[15487]= -2063024031;
assign addr[15488]= -2040479063;
assign addr[15489]= -2015345591;
assign addr[15490]= -1987655498;
assign addr[15491]= -1957443913;
assign addr[15492]= -1924749160;
assign addr[15493]= -1889612716;
assign addr[15494]= -1852079154;
assign addr[15495]= -1812196087;
assign addr[15496]= -1770014111;
assign addr[15497]= -1725586737;
assign addr[15498]= -1678970324;
assign addr[15499]= -1630224009;
assign addr[15500]= -1579409630;
assign addr[15501]= -1526591649;
assign addr[15502]= -1471837070;
assign addr[15503]= -1415215352;
assign addr[15504]= -1356798326;
assign addr[15505]= -1296660098;
assign addr[15506]= -1234876957;
assign addr[15507]= -1171527280;
assign addr[15508]= -1106691431;
assign addr[15509]= -1040451659;
assign addr[15510]= -972891995;
assign addr[15511]= -904098143;
assign addr[15512]= -834157373;
assign addr[15513]= -763158411;
assign addr[15514]= -691191324;
assign addr[15515]= -618347408;
assign addr[15516]= -544719071;
assign addr[15517]= -470399716;
assign addr[15518]= -395483624;
assign addr[15519]= -320065829;
assign addr[15520]= -244242007;
assign addr[15521]= -168108346;
assign addr[15522]= -91761426;
assign addr[15523]= -15298099;
assign addr[15524]= 61184634;
assign addr[15525]= 137589750;
assign addr[15526]= 213820322;
assign addr[15527]= 289779648;
assign addr[15528]= 365371365;
assign addr[15529]= 440499581;
assign addr[15530]= 515068990;
assign addr[15531]= 588984994;
assign addr[15532]= 662153826;
assign addr[15533]= 734482665;
assign addr[15534]= 805879757;
assign addr[15535]= 876254528;
assign addr[15536]= 945517704;
assign addr[15537]= 1013581418;
assign addr[15538]= 1080359326;
assign addr[15539]= 1145766716;
assign addr[15540]= 1209720613;
assign addr[15541]= 1272139887;
assign addr[15542]= 1332945355;
assign addr[15543]= 1392059879;
assign addr[15544]= 1449408469;
assign addr[15545]= 1504918373;
assign addr[15546]= 1558519173;
assign addr[15547]= 1610142873;
assign addr[15548]= 1659723983;
assign addr[15549]= 1707199606;
assign addr[15550]= 1752509516;
assign addr[15551]= 1795596234;
assign addr[15552]= 1836405100;
assign addr[15553]= 1874884346;
assign addr[15554]= 1910985158;
assign addr[15555]= 1944661739;
assign addr[15556]= 1975871368;
assign addr[15557]= 2004574453;
assign addr[15558]= 2030734582;
assign addr[15559]= 2054318569;
assign addr[15560]= 2075296495;
assign addr[15561]= 2093641749;
assign addr[15562]= 2109331059;
assign addr[15563]= 2122344521;
assign addr[15564]= 2132665626;
assign addr[15565]= 2140281282;
assign addr[15566]= 2145181827;
assign addr[15567]= 2147361045;
assign addr[15568]= 2146816171;
assign addr[15569]= 2143547897;
assign addr[15570]= 2137560369;
assign addr[15571]= 2128861181;
assign addr[15572]= 2117461370;
assign addr[15573]= 2103375398;
assign addr[15574]= 2086621133;
assign addr[15575]= 2067219829;
assign addr[15576]= 2045196100;
assign addr[15577]= 2020577882;
assign addr[15578]= 1993396407;
assign addr[15579]= 1963686155;
assign addr[15580]= 1931484818;
assign addr[15581]= 1896833245;
assign addr[15582]= 1859775393;
assign addr[15583]= 1820358275;
assign addr[15584]= 1778631892;
assign addr[15585]= 1734649179;
assign addr[15586]= 1688465931;
assign addr[15587]= 1640140734;
assign addr[15588]= 1589734894;
assign addr[15589]= 1537312353;
assign addr[15590]= 1482939614;
assign addr[15591]= 1426685652;
assign addr[15592]= 1368621831;
assign addr[15593]= 1308821808;
assign addr[15594]= 1247361445;
assign addr[15595]= 1184318708;
assign addr[15596]= 1119773573;
assign addr[15597]= 1053807919;
assign addr[15598]= 986505429;
assign addr[15599]= 917951481;
assign addr[15600]= 848233042;
assign addr[15601]= 777438554;
assign addr[15602]= 705657826;
assign addr[15603]= 632981917;
assign addr[15604]= 559503022;
assign addr[15605]= 485314355;
assign addr[15606]= 410510029;
assign addr[15607]= 335184940;
assign addr[15608]= 259434643;
assign addr[15609]= 183355234;
assign addr[15610]= 107043224;
assign addr[15611]= 30595422;
assign addr[15612]= -45891193;
assign addr[15613]= -122319591;
assign addr[15614]= -198592817;
assign addr[15615]= -274614114;
assign addr[15616]= -350287041;
assign addr[15617]= -425515602;
assign addr[15618]= -500204365;
assign addr[15619]= -574258580;
assign addr[15620]= -647584304;
assign addr[15621]= -720088517;
assign addr[15622]= -791679244;
assign addr[15623]= -862265664;
assign addr[15624]= -931758235;
assign addr[15625]= -1000068799;
assign addr[15626]= -1067110699;
assign addr[15627]= -1132798888;
assign addr[15628]= -1197050035;
assign addr[15629]= -1259782632;
assign addr[15630]= -1320917099;
assign addr[15631]= -1380375881;
assign addr[15632]= -1438083551;
assign addr[15633]= -1493966902;
assign addr[15634]= -1547955041;
assign addr[15635]= -1599979481;
assign addr[15636]= -1649974225;
assign addr[15637]= -1697875851;
assign addr[15638]= -1743623590;
assign addr[15639]= -1787159411;
assign addr[15640]= -1828428082;
assign addr[15641]= -1867377253;
assign addr[15642]= -1903957513;
assign addr[15643]= -1938122457;
assign addr[15644]= -1969828744;
assign addr[15645]= -1999036154;
assign addr[15646]= -2025707632;
assign addr[15647]= -2049809346;
assign addr[15648]= -2071310720;
assign addr[15649]= -2090184478;
assign addr[15650]= -2106406677;
assign addr[15651]= -2119956737;
assign addr[15652]= -2130817471;
assign addr[15653]= -2138975100;
assign addr[15654]= -2144419275;
assign addr[15655]= -2147143090;
assign addr[15656]= -2147143090;
assign addr[15657]= -2144419275;
assign addr[15658]= -2138975100;
assign addr[15659]= -2130817471;
assign addr[15660]= -2119956737;
assign addr[15661]= -2106406677;
assign addr[15662]= -2090184478;
assign addr[15663]= -2071310720;
assign addr[15664]= -2049809346;
assign addr[15665]= -2025707632;
assign addr[15666]= -1999036154;
assign addr[15667]= -1969828744;
assign addr[15668]= -1938122457;
assign addr[15669]= -1903957513;
assign addr[15670]= -1867377253;
assign addr[15671]= -1828428082;
assign addr[15672]= -1787159411;
assign addr[15673]= -1743623590;
assign addr[15674]= -1697875851;
assign addr[15675]= -1649974225;
assign addr[15676]= -1599979481;
assign addr[15677]= -1547955041;
assign addr[15678]= -1493966902;
assign addr[15679]= -1438083551;
assign addr[15680]= -1380375881;
assign addr[15681]= -1320917099;
assign addr[15682]= -1259782632;
assign addr[15683]= -1197050035;
assign addr[15684]= -1132798888;
assign addr[15685]= -1067110699;
assign addr[15686]= -1000068799;
assign addr[15687]= -931758235;
assign addr[15688]= -862265664;
assign addr[15689]= -791679244;
assign addr[15690]= -720088517;
assign addr[15691]= -647584304;
assign addr[15692]= -574258580;
assign addr[15693]= -500204365;
assign addr[15694]= -425515602;
assign addr[15695]= -350287041;
assign addr[15696]= -274614114;
assign addr[15697]= -198592817;
assign addr[15698]= -122319591;
assign addr[15699]= -45891193;
assign addr[15700]= 30595422;
assign addr[15701]= 107043224;
assign addr[15702]= 183355234;
assign addr[15703]= 259434643;
assign addr[15704]= 335184940;
assign addr[15705]= 410510029;
assign addr[15706]= 485314355;
assign addr[15707]= 559503022;
assign addr[15708]= 632981917;
assign addr[15709]= 705657826;
assign addr[15710]= 777438554;
assign addr[15711]= 848233042;
assign addr[15712]= 917951481;
assign addr[15713]= 986505429;
assign addr[15714]= 1053807919;
assign addr[15715]= 1119773573;
assign addr[15716]= 1184318708;
assign addr[15717]= 1247361445;
assign addr[15718]= 1308821808;
assign addr[15719]= 1368621831;
assign addr[15720]= 1426685652;
assign addr[15721]= 1482939614;
assign addr[15722]= 1537312353;
assign addr[15723]= 1589734894;
assign addr[15724]= 1640140734;
assign addr[15725]= 1688465931;
assign addr[15726]= 1734649179;
assign addr[15727]= 1778631892;
assign addr[15728]= 1820358275;
assign addr[15729]= 1859775393;
assign addr[15730]= 1896833245;
assign addr[15731]= 1931484818;
assign addr[15732]= 1963686155;
assign addr[15733]= 1993396407;
assign addr[15734]= 2020577882;
assign addr[15735]= 2045196100;
assign addr[15736]= 2067219829;
assign addr[15737]= 2086621133;
assign addr[15738]= 2103375398;
assign addr[15739]= 2117461370;
assign addr[15740]= 2128861181;
assign addr[15741]= 2137560369;
assign addr[15742]= 2143547897;
assign addr[15743]= 2146816171;
assign addr[15744]= 2147361045;
assign addr[15745]= 2145181827;
assign addr[15746]= 2140281282;
assign addr[15747]= 2132665626;
assign addr[15748]= 2122344521;
assign addr[15749]= 2109331059;
assign addr[15750]= 2093641749;
assign addr[15751]= 2075296495;
assign addr[15752]= 2054318569;
assign addr[15753]= 2030734582;
assign addr[15754]= 2004574453;
assign addr[15755]= 1975871368;
assign addr[15756]= 1944661739;
assign addr[15757]= 1910985158;
assign addr[15758]= 1874884346;
assign addr[15759]= 1836405100;
assign addr[15760]= 1795596234;
assign addr[15761]= 1752509516;
assign addr[15762]= 1707199606;
assign addr[15763]= 1659723983;
assign addr[15764]= 1610142873;
assign addr[15765]= 1558519173;
assign addr[15766]= 1504918373;
assign addr[15767]= 1449408469;
assign addr[15768]= 1392059879;
assign addr[15769]= 1332945355;
assign addr[15770]= 1272139887;
assign addr[15771]= 1209720613;
assign addr[15772]= 1145766716;
assign addr[15773]= 1080359326;
assign addr[15774]= 1013581418;
assign addr[15775]= 945517704;
assign addr[15776]= 876254528;
assign addr[15777]= 805879757;
assign addr[15778]= 734482665;
assign addr[15779]= 662153826;
assign addr[15780]= 588984994;
assign addr[15781]= 515068990;
assign addr[15782]= 440499581;
assign addr[15783]= 365371365;
assign addr[15784]= 289779648;
assign addr[15785]= 213820322;
assign addr[15786]= 137589750;
assign addr[15787]= 61184634;
assign addr[15788]= -15298099;
assign addr[15789]= -91761426;
assign addr[15790]= -168108346;
assign addr[15791]= -244242007;
assign addr[15792]= -320065829;
assign addr[15793]= -395483624;
assign addr[15794]= -470399716;
assign addr[15795]= -544719071;
assign addr[15796]= -618347408;
assign addr[15797]= -691191324;
assign addr[15798]= -763158411;
assign addr[15799]= -834157373;
assign addr[15800]= -904098143;
assign addr[15801]= -972891995;
assign addr[15802]= -1040451659;
assign addr[15803]= -1106691431;
assign addr[15804]= -1171527280;
assign addr[15805]= -1234876957;
assign addr[15806]= -1296660098;
assign addr[15807]= -1356798326;
assign addr[15808]= -1415215352;
assign addr[15809]= -1471837070;
assign addr[15810]= -1526591649;
assign addr[15811]= -1579409630;
assign addr[15812]= -1630224009;
assign addr[15813]= -1678970324;
assign addr[15814]= -1725586737;
assign addr[15815]= -1770014111;
assign addr[15816]= -1812196087;
assign addr[15817]= -1852079154;
assign addr[15818]= -1889612716;
assign addr[15819]= -1924749160;
assign addr[15820]= -1957443913;
assign addr[15821]= -1987655498;
assign addr[15822]= -2015345591;
assign addr[15823]= -2040479063;
assign addr[15824]= -2063024031;
assign addr[15825]= -2082951896;
assign addr[15826]= -2100237377;
assign addr[15827]= -2114858546;
assign addr[15828]= -2126796855;
assign addr[15829]= -2136037160;
assign addr[15830]= -2142567738;
assign addr[15831]= -2146380306;
assign addr[15832]= -2147470025;
assign addr[15833]= -2145835515;
assign addr[15834]= -2141478848;
assign addr[15835]= -2134405552;
assign addr[15836]= -2124624598;
assign addr[15837]= -2112148396;
assign addr[15838]= -2096992772;
assign addr[15839]= -2079176953;
assign addr[15840]= -2058723538;
assign addr[15841]= -2035658475;
assign addr[15842]= -2010011024;
assign addr[15843]= -1981813720;
assign addr[15844]= -1951102334;
assign addr[15845]= -1917915825;
assign addr[15846]= -1882296293;
assign addr[15847]= -1844288924;
assign addr[15848]= -1803941934;
assign addr[15849]= -1761306505;
assign addr[15850]= -1716436725;
assign addr[15851]= -1669389513;
assign addr[15852]= -1620224553;
assign addr[15853]= -1569004214;
assign addr[15854]= -1515793473;
assign addr[15855]= -1460659832;
assign addr[15856]= -1403673233;
assign addr[15857]= -1344905966;
assign addr[15858]= -1284432584;
assign addr[15859]= -1222329801;
assign addr[15860]= -1158676398;
assign addr[15861]= -1093553126;
assign addr[15862]= -1027042599;
assign addr[15863]= -959229189;
assign addr[15864]= -890198924;
assign addr[15865]= -820039373;
assign addr[15866]= -748839539;
assign addr[15867]= -676689746;
assign addr[15868]= -603681519;
assign addr[15869]= -529907477;
assign addr[15870]= -455461206;
assign addr[15871]= -380437148;
assign addr[15872]= -304930476;
assign addr[15873]= -229036977;
assign addr[15874]= -152852926;
assign addr[15875]= -76474970;
assign addr[15876]= 0;
assign addr[15877]= 76474970;
assign addr[15878]= 152852926;
assign addr[15879]= 229036977;
assign addr[15880]= 304930476;
assign addr[15881]= 380437148;
assign addr[15882]= 455461206;
assign addr[15883]= 529907477;
assign addr[15884]= 603681519;
assign addr[15885]= 676689746;
assign addr[15886]= 748839539;
assign addr[15887]= 820039373;
assign addr[15888]= 890198924;
assign addr[15889]= 959229189;
assign addr[15890]= 1027042599;
assign addr[15891]= 1093553126;
assign addr[15892]= 1158676398;
assign addr[15893]= 1222329801;
assign addr[15894]= 1284432584;
assign addr[15895]= 1344905966;
assign addr[15896]= 1403673233;
assign addr[15897]= 1460659832;
assign addr[15898]= 1515793473;
assign addr[15899]= 1569004214;
assign addr[15900]= 1620224553;
assign addr[15901]= 1669389513;
assign addr[15902]= 1716436725;
assign addr[15903]= 1761306505;
assign addr[15904]= 1803941934;
assign addr[15905]= 1844288924;
assign addr[15906]= 1882296293;
assign addr[15907]= 1917915825;
assign addr[15908]= 1951102334;
assign addr[15909]= 1981813720;
assign addr[15910]= 2010011024;
assign addr[15911]= 2035658475;
assign addr[15912]= 2058723538;
assign addr[15913]= 2079176953;
assign addr[15914]= 2096992772;
assign addr[15915]= 2112148396;
assign addr[15916]= 2124624598;
assign addr[15917]= 2134405552;
assign addr[15918]= 2141478848;
assign addr[15919]= 2145835515;
assign addr[15920]= 2147470025;
assign addr[15921]= 2146380306;
assign addr[15922]= 2142567738;
assign addr[15923]= 2136037160;
assign addr[15924]= 2126796855;
assign addr[15925]= 2114858546;
assign addr[15926]= 2100237377;
assign addr[15927]= 2082951896;
assign addr[15928]= 2063024031;
assign addr[15929]= 2040479063;
assign addr[15930]= 2015345591;
assign addr[15931]= 1987655498;
assign addr[15932]= 1957443913;
assign addr[15933]= 1924749160;
assign addr[15934]= 1889612716;
assign addr[15935]= 1852079154;
assign addr[15936]= 1812196087;
assign addr[15937]= 1770014111;
assign addr[15938]= 1725586737;
assign addr[15939]= 1678970324;
assign addr[15940]= 1630224009;
assign addr[15941]= 1579409630;
assign addr[15942]= 1526591649;
assign addr[15943]= 1471837070;
assign addr[15944]= 1415215352;
assign addr[15945]= 1356798326;
assign addr[15946]= 1296660098;
assign addr[15947]= 1234876957;
assign addr[15948]= 1171527280;
assign addr[15949]= 1106691431;
assign addr[15950]= 1040451659;
assign addr[15951]= 972891995;
assign addr[15952]= 904098143;
assign addr[15953]= 834157373;
assign addr[15954]= 763158411;
assign addr[15955]= 691191324;
assign addr[15956]= 618347408;
assign addr[15957]= 544719071;
assign addr[15958]= 470399716;
assign addr[15959]= 395483624;
assign addr[15960]= 320065829;
assign addr[15961]= 244242007;
assign addr[15962]= 168108346;
assign addr[15963]= 91761426;
assign addr[15964]= 15298099;
assign addr[15965]= -61184634;
assign addr[15966]= -137589750;
assign addr[15967]= -213820322;
assign addr[15968]= -289779648;
assign addr[15969]= -365371365;
assign addr[15970]= -440499581;
assign addr[15971]= -515068990;
assign addr[15972]= -588984994;
assign addr[15973]= -662153826;
assign addr[15974]= -734482665;
assign addr[15975]= -805879757;
assign addr[15976]= -876254528;
assign addr[15977]= -945517704;
assign addr[15978]= -1013581418;
assign addr[15979]= -1080359326;
assign addr[15980]= -1145766716;
assign addr[15981]= -1209720613;
assign addr[15982]= -1272139887;
assign addr[15983]= -1332945355;
assign addr[15984]= -1392059879;
assign addr[15985]= -1449408469;
assign addr[15986]= -1504918373;
assign addr[15987]= -1558519173;
assign addr[15988]= -1610142873;
assign addr[15989]= -1659723983;
assign addr[15990]= -1707199606;
assign addr[15991]= -1752509516;
assign addr[15992]= -1795596234;
assign addr[15993]= -1836405100;
assign addr[15994]= -1874884346;
assign addr[15995]= -1910985158;
assign addr[15996]= -1944661739;
assign addr[15997]= -1975871368;
assign addr[15998]= -2004574453;
assign addr[15999]= -2030734582;
assign addr[16000]= -2054318569;
assign addr[16001]= -2075296495;
assign addr[16002]= -2093641749;
assign addr[16003]= -2109331059;
assign addr[16004]= -2122344521;
assign addr[16005]= -2132665626;
assign addr[16006]= -2140281282;
assign addr[16007]= -2145181827;
assign addr[16008]= -2147361045;
assign addr[16009]= -2146816171;
assign addr[16010]= -2143547897;
assign addr[16011]= -2137560369;
assign addr[16012]= -2128861181;
assign addr[16013]= -2117461370;
assign addr[16014]= -2103375398;
assign addr[16015]= -2086621133;
assign addr[16016]= -2067219829;
assign addr[16017]= -2045196100;
assign addr[16018]= -2020577882;
assign addr[16019]= -1993396407;
assign addr[16020]= -1963686155;
assign addr[16021]= -1931484818;
assign addr[16022]= -1896833245;
assign addr[16023]= -1859775393;
assign addr[16024]= -1820358275;
assign addr[16025]= -1778631892;
assign addr[16026]= -1734649179;
assign addr[16027]= -1688465931;
assign addr[16028]= -1640140734;
assign addr[16029]= -1589734894;
assign addr[16030]= -1537312353;
assign addr[16031]= -1482939614;
assign addr[16032]= -1426685652;
assign addr[16033]= -1368621831;
assign addr[16034]= -1308821808;
assign addr[16035]= -1247361445;
assign addr[16036]= -1184318708;
assign addr[16037]= -1119773573;
assign addr[16038]= -1053807919;
assign addr[16039]= -986505429;
assign addr[16040]= -917951481;
assign addr[16041]= -848233042;
assign addr[16042]= -777438554;
assign addr[16043]= -705657826;
assign addr[16044]= -632981917;
assign addr[16045]= -559503022;
assign addr[16046]= -485314355;
assign addr[16047]= -410510029;
assign addr[16048]= -335184940;
assign addr[16049]= -259434643;
assign addr[16050]= -183355234;
assign addr[16051]= -107043224;
assign addr[16052]= -30595422;
assign addr[16053]= 45891193;
assign addr[16054]= 122319591;
assign addr[16055]= 198592817;
assign addr[16056]= 274614114;
assign addr[16057]= 350287041;
assign addr[16058]= 425515602;
assign addr[16059]= 500204365;
assign addr[16060]= 574258580;
assign addr[16061]= 647584304;
assign addr[16062]= 720088517;
assign addr[16063]= 791679244;
assign addr[16064]= 862265664;
assign addr[16065]= 931758235;
assign addr[16066]= 1000068799;
assign addr[16067]= 1067110699;
assign addr[16068]= 1132798888;
assign addr[16069]= 1197050035;
assign addr[16070]= 1259782632;
assign addr[16071]= 1320917099;
assign addr[16072]= 1380375881;
assign addr[16073]= 1438083551;
assign addr[16074]= 1493966902;
assign addr[16075]= 1547955041;
assign addr[16076]= 1599979481;
assign addr[16077]= 1649974225;
assign addr[16078]= 1697875851;
assign addr[16079]= 1743623590;
assign addr[16080]= 1787159411;
assign addr[16081]= 1828428082;
assign addr[16082]= 1867377253;
assign addr[16083]= 1903957513;
assign addr[16084]= 1938122457;
assign addr[16085]= 1969828744;
assign addr[16086]= 1999036154;
assign addr[16087]= 2025707632;
assign addr[16088]= 2049809346;
assign addr[16089]= 2071310720;
assign addr[16090]= 2090184478;
assign addr[16091]= 2106406677;
assign addr[16092]= 2119956737;
assign addr[16093]= 2130817471;
assign addr[16094]= 2138975100;
assign addr[16095]= 2144419275;
assign addr[16096]= 2147143090;
assign addr[16097]= 2147143090;
assign addr[16098]= 2144419275;
assign addr[16099]= 2138975100;
assign addr[16100]= 2130817471;
assign addr[16101]= 2119956737;
assign addr[16102]= 2106406677;
assign addr[16103]= 2090184478;
assign addr[16104]= 2071310720;
assign addr[16105]= 2049809346;
assign addr[16106]= 2025707632;
assign addr[16107]= 1999036154;
assign addr[16108]= 1969828744;
assign addr[16109]= 1938122457;
assign addr[16110]= 1903957513;
assign addr[16111]= 1867377253;
assign addr[16112]= 1828428082;
assign addr[16113]= 1787159411;
assign addr[16114]= 1743623590;
assign addr[16115]= 1697875851;
assign addr[16116]= 1649974225;
assign addr[16117]= 1599979481;
assign addr[16118]= 1547955041;
assign addr[16119]= 1493966902;
assign addr[16120]= 1438083551;
assign addr[16121]= 1380375881;
assign addr[16122]= 1320917099;
assign addr[16123]= 1259782632;
assign addr[16124]= 1197050035;
assign addr[16125]= 1132798888;
assign addr[16126]= 1067110699;
assign addr[16127]= 1000068799;
assign addr[16128]= 931758235;
assign addr[16129]= 862265664;
assign addr[16130]= 791679244;
assign addr[16131]= 720088517;
assign addr[16132]= 647584304;
assign addr[16133]= 574258580;
assign addr[16134]= 500204365;
assign addr[16135]= 425515602;
assign addr[16136]= 350287041;
assign addr[16137]= 274614114;
assign addr[16138]= 198592817;
assign addr[16139]= 122319591;
assign addr[16140]= 45891193;
assign addr[16141]= -30595422;
assign addr[16142]= -107043224;
assign addr[16143]= -183355234;
assign addr[16144]= -259434643;
assign addr[16145]= -335184940;
assign addr[16146]= -410510029;
assign addr[16147]= -485314355;
assign addr[16148]= -559503022;
assign addr[16149]= -632981917;
assign addr[16150]= -705657826;
assign addr[16151]= -777438554;
assign addr[16152]= -848233042;
assign addr[16153]= -917951481;
assign addr[16154]= -986505429;
assign addr[16155]= -1053807919;
assign addr[16156]= -1119773573;
assign addr[16157]= -1184318708;
assign addr[16158]= -1247361445;
assign addr[16159]= -1308821808;
assign addr[16160]= -1368621831;
assign addr[16161]= -1426685652;
assign addr[16162]= -1482939614;
assign addr[16163]= -1537312353;
assign addr[16164]= -1589734894;
assign addr[16165]= -1640140734;
assign addr[16166]= -1688465931;
assign addr[16167]= -1734649179;
assign addr[16168]= -1778631892;
assign addr[16169]= -1820358275;
assign addr[16170]= -1859775393;
assign addr[16171]= -1896833245;
assign addr[16172]= -1931484818;
assign addr[16173]= -1963686155;
assign addr[16174]= -1993396407;
assign addr[16175]= -2020577882;
assign addr[16176]= -2045196100;
assign addr[16177]= -2067219829;
assign addr[16178]= -2086621133;
assign addr[16179]= -2103375398;
assign addr[16180]= -2117461370;
assign addr[16181]= -2128861181;
assign addr[16182]= -2137560369;
assign addr[16183]= -2143547897;
assign addr[16184]= -2146816171;
assign addr[16185]= -2147361045;
assign addr[16186]= -2145181827;
assign addr[16187]= -2140281282;
assign addr[16188]= -2132665626;
assign addr[16189]= -2122344521;
assign addr[16190]= -2109331059;
assign addr[16191]= -2093641749;
assign addr[16192]= -2075296495;
assign addr[16193]= -2054318569;
assign addr[16194]= -2030734582;
assign addr[16195]= -2004574453;
assign addr[16196]= -1975871368;
assign addr[16197]= -1944661739;
assign addr[16198]= -1910985158;
assign addr[16199]= -1874884346;
assign addr[16200]= -1836405100;
assign addr[16201]= -1795596234;
assign addr[16202]= -1752509516;
assign addr[16203]= -1707199606;
assign addr[16204]= -1659723983;
assign addr[16205]= -1610142873;
assign addr[16206]= -1558519173;
assign addr[16207]= -1504918373;
assign addr[16208]= -1449408469;
assign addr[16209]= -1392059879;
assign addr[16210]= -1332945355;
assign addr[16211]= -1272139887;
assign addr[16212]= -1209720613;
assign addr[16213]= -1145766716;
assign addr[16214]= -1080359326;
assign addr[16215]= -1013581418;
assign addr[16216]= -945517704;
assign addr[16217]= -876254528;
assign addr[16218]= -805879757;
assign addr[16219]= -734482665;
assign addr[16220]= -662153826;
assign addr[16221]= -588984994;
assign addr[16222]= -515068990;
assign addr[16223]= -440499581;
assign addr[16224]= -365371365;
assign addr[16225]= -289779648;
assign addr[16226]= -213820322;
assign addr[16227]= -137589750;
assign addr[16228]= -61184634;
assign addr[16229]= 15298099;
assign addr[16230]= 91761426;
assign addr[16231]= 168108346;
assign addr[16232]= 244242007;
assign addr[16233]= 320065829;
assign addr[16234]= 395483624;
assign addr[16235]= 470399716;
assign addr[16236]= 544719071;
assign addr[16237]= 618347408;
assign addr[16238]= 691191324;
assign addr[16239]= 763158411;
assign addr[16240]= 834157373;
assign addr[16241]= 904098143;
assign addr[16242]= 972891995;
assign addr[16243]= 1040451659;
assign addr[16244]= 1106691431;
assign addr[16245]= 1171527280;
assign addr[16246]= 1234876957;
assign addr[16247]= 1296660098;
assign addr[16248]= 1356798326;
assign addr[16249]= 1415215352;
assign addr[16250]= 1471837070;
assign addr[16251]= 1526591649;
assign addr[16252]= 1579409630;
assign addr[16253]= 1630224009;
assign addr[16254]= 1678970324;
assign addr[16255]= 1725586737;
assign addr[16256]= 1770014111;
assign addr[16257]= 1812196087;
assign addr[16258]= 1852079154;
assign addr[16259]= 1889612716;
assign addr[16260]= 1924749160;
assign addr[16261]= 1957443913;
assign addr[16262]= 1987655498;
assign addr[16263]= 2015345591;
assign addr[16264]= 2040479063;
assign addr[16265]= 2063024031;
assign addr[16266]= 2082951896;
assign addr[16267]= 2100237377;
assign addr[16268]= 2114858546;
assign addr[16269]= 2126796855;
assign addr[16270]= 2136037160;
assign addr[16271]= 2142567738;
assign addr[16272]= 2146380306;
assign addr[16273]= 2147470025;
assign addr[16274]= 2145835515;
assign addr[16275]= 2141478848;
assign addr[16276]= 2134405552;
assign addr[16277]= 2124624598;
assign addr[16278]= 2112148396;
assign addr[16279]= 2096992772;
assign addr[16280]= 2079176953;
assign addr[16281]= 2058723538;
assign addr[16282]= 2035658475;
assign addr[16283]= 2010011024;
assign addr[16284]= 1981813720;
assign addr[16285]= 1951102334;
assign addr[16286]= 1917915825;
assign addr[16287]= 1882296293;
assign addr[16288]= 1844288924;
assign addr[16289]= 1803941934;
assign addr[16290]= 1761306505;
assign addr[16291]= 1716436725;
assign addr[16292]= 1669389513;
assign addr[16293]= 1620224553;
assign addr[16294]= 1569004214;
assign addr[16295]= 1515793473;
assign addr[16296]= 1460659832;
assign addr[16297]= 1403673233;
assign addr[16298]= 1344905966;
assign addr[16299]= 1284432584;
assign addr[16300]= 1222329801;
assign addr[16301]= 1158676398;
assign addr[16302]= 1093553126;
assign addr[16303]= 1027042599;
assign addr[16304]= 959229189;
assign addr[16305]= 890198924;
assign addr[16306]= 820039373;
assign addr[16307]= 748839539;
assign addr[16308]= 676689746;
assign addr[16309]= 603681519;
assign addr[16310]= 529907477;
assign addr[16311]= 455461206;
assign addr[16312]= 380437148;
assign addr[16313]= 304930476;
assign addr[16314]= 229036977;
assign addr[16315]= 152852926;
assign addr[16316]= 76474970;
assign addr[16317]= 0;
assign addr[16318]= -76474970;
assign addr[16319]= -152852926;
assign addr[16320]= -229036977;
assign addr[16321]= -304930476;
assign addr[16322]= -380437148;
assign addr[16323]= -455461206;
assign addr[16324]= -529907477;
assign addr[16325]= -603681519;
assign addr[16326]= -676689746;
assign addr[16327]= -748839539;
assign addr[16328]= -820039373;
assign addr[16329]= -890198924;
assign addr[16330]= -959229189;
assign addr[16331]= -1027042599;
assign addr[16332]= -1093553126;
assign addr[16333]= -1158676398;
assign addr[16334]= -1222329801;
assign addr[16335]= -1284432584;
assign addr[16336]= -1344905966;
assign addr[16337]= -1403673233;
assign addr[16338]= -1460659832;
assign addr[16339]= -1515793473;
assign addr[16340]= -1569004214;
assign addr[16341]= -1620224553;
assign addr[16342]= -1669389513;
assign addr[16343]= -1716436725;
assign addr[16344]= -1761306505;
assign addr[16345]= -1803941934;
assign addr[16346]= -1844288924;
assign addr[16347]= -1882296293;
assign addr[16348]= -1917915825;
assign addr[16349]= -1951102334;
assign addr[16350]= -1981813720;
assign addr[16351]= -2010011024;
assign addr[16352]= -2035658475;
assign addr[16353]= -2058723538;
assign addr[16354]= -2079176953;
assign addr[16355]= -2096992772;
assign addr[16356]= -2112148396;
assign addr[16357]= -2124624598;
assign addr[16358]= -2134405552;
assign addr[16359]= -2141478848;
assign addr[16360]= -2145835515;
assign addr[16361]= -2147470025;
assign addr[16362]= -2146380306;
assign addr[16363]= -2142567738;
assign addr[16364]= -2136037160;
assign addr[16365]= -2126796855;
assign addr[16366]= -2114858546;
assign addr[16367]= -2100237377;
assign addr[16368]= -2082951896;
assign addr[16369]= -2063024031;
assign addr[16370]= -2040479063;
assign addr[16371]= -2015345591;
assign addr[16372]= -1987655498;
assign addr[16373]= -1957443913;
assign addr[16374]= -1924749160;
assign addr[16375]= -1889612716;
assign addr[16376]= -1852079154;
assign addr[16377]= -1812196087;
assign addr[16378]= -1770014111;
assign addr[16379]= -1725586737;
assign addr[16380]= -1678970324;
assign addr[16381]= -1630224009;
assign addr[16382]= -1579409630;
assign addr[16383]= -1526591649;
assign addr[16384]= -1471837070;
assign addr[16385]= -1415215352;
assign addr[16386]= -1356798326;
assign addr[16387]= -1296660098;
assign addr[16388]= -1234876957;
assign addr[16389]= -1171527280;
assign addr[16390]= -1106691431;
assign addr[16391]= -1040451659;
assign addr[16392]= -972891995;
assign addr[16393]= -904098143;
assign addr[16394]= -834157373;
assign addr[16395]= -763158411;
assign addr[16396]= -691191324;
assign addr[16397]= -618347408;
assign addr[16398]= -544719071;
assign addr[16399]= -470399716;
assign addr[16400]= -395483624;
assign addr[16401]= -320065829;
assign addr[16402]= -244242007;
assign addr[16403]= -168108346;
assign addr[16404]= -91761426;
assign addr[16405]= -15298099;
assign addr[16406]= 61184634;
assign addr[16407]= 137589750;
assign addr[16408]= 213820322;
assign addr[16409]= 289779648;
assign addr[16410]= 365371365;
assign addr[16411]= 440499581;
assign addr[16412]= 515068990;
assign addr[16413]= 588984994;
assign addr[16414]= 662153826;
assign addr[16415]= 734482665;
assign addr[16416]= 805879757;
assign addr[16417]= 876254528;
assign addr[16418]= 945517704;
assign addr[16419]= 1013581418;
assign addr[16420]= 1080359326;
assign addr[16421]= 1145766716;
assign addr[16422]= 1209720613;
assign addr[16423]= 1272139887;
assign addr[16424]= 1332945355;
assign addr[16425]= 1392059879;
assign addr[16426]= 1449408469;
assign addr[16427]= 1504918373;
assign addr[16428]= 1558519173;
assign addr[16429]= 1610142873;
assign addr[16430]= 1659723983;
assign addr[16431]= 1707199606;
assign addr[16432]= 1752509516;
assign addr[16433]= 1795596234;
assign addr[16434]= 1836405100;
assign addr[16435]= 1874884346;
assign addr[16436]= 1910985158;
assign addr[16437]= 1944661739;
assign addr[16438]= 1975871368;
assign addr[16439]= 2004574453;
assign addr[16440]= 2030734582;
assign addr[16441]= 2054318569;
assign addr[16442]= 2075296495;
assign addr[16443]= 2093641749;
assign addr[16444]= 2109331059;
assign addr[16445]= 2122344521;
assign addr[16446]= 2132665626;
assign addr[16447]= 2140281282;
assign addr[16448]= 2145181827;
assign addr[16449]= 2147361045;
assign addr[16450]= 2146816171;
assign addr[16451]= 2143547897;
assign addr[16452]= 2137560369;
assign addr[16453]= 2128861181;
assign addr[16454]= 2117461370;
assign addr[16455]= 2103375398;
assign addr[16456]= 2086621133;
assign addr[16457]= 2067219829;
assign addr[16458]= 2045196100;
assign addr[16459]= 2020577882;
assign addr[16460]= 1993396407;
assign addr[16461]= 1963686155;
assign addr[16462]= 1931484818;
assign addr[16463]= 1896833245;
assign addr[16464]= 1859775393;
assign addr[16465]= 1820358275;
assign addr[16466]= 1778631892;
assign addr[16467]= 1734649179;
assign addr[16468]= 1688465931;
assign addr[16469]= 1640140734;
assign addr[16470]= 1589734894;
assign addr[16471]= 1537312353;
assign addr[16472]= 1482939614;
assign addr[16473]= 1426685652;
assign addr[16474]= 1368621831;
assign addr[16475]= 1308821808;
assign addr[16476]= 1247361445;
assign addr[16477]= 1184318708;
assign addr[16478]= 1119773573;
assign addr[16479]= 1053807919;
assign addr[16480]= 986505429;
assign addr[16481]= 917951481;
assign addr[16482]= 848233042;
assign addr[16483]= 777438554;
assign addr[16484]= 705657826;
assign addr[16485]= 632981917;
assign addr[16486]= 559503022;
assign addr[16487]= 485314355;
assign addr[16488]= 410510029;
assign addr[16489]= 335184940;
assign addr[16490]= 259434643;
assign addr[16491]= 183355234;
assign addr[16492]= 107043224;
assign addr[16493]= 30595422;
assign addr[16494]= -45891193;
assign addr[16495]= -122319591;
assign addr[16496]= -198592817;
assign addr[16497]= -274614114;
assign addr[16498]= -350287041;
assign addr[16499]= -425515602;
assign addr[16500]= -500204365;
assign addr[16501]= -574258580;
assign addr[16502]= -647584304;
assign addr[16503]= -720088517;
assign addr[16504]= -791679244;
assign addr[16505]= -862265664;
assign addr[16506]= -931758235;
assign addr[16507]= -1000068799;
assign addr[16508]= -1067110699;
assign addr[16509]= -1132798888;
assign addr[16510]= -1197050035;
assign addr[16511]= -1259782632;
assign addr[16512]= -1320917099;
assign addr[16513]= -1380375881;
assign addr[16514]= -1438083551;
assign addr[16515]= -1493966902;
assign addr[16516]= -1547955041;
assign addr[16517]= -1599979481;
assign addr[16518]= -1649974225;
assign addr[16519]= -1697875851;
assign addr[16520]= -1743623590;
assign addr[16521]= -1787159411;
assign addr[16522]= -1828428082;
assign addr[16523]= -1867377253;
assign addr[16524]= -1903957513;
assign addr[16525]= -1938122457;
assign addr[16526]= -1969828744;
assign addr[16527]= -1999036154;
assign addr[16528]= -2025707632;
assign addr[16529]= -2049809346;
assign addr[16530]= -2071310720;
assign addr[16531]= -2090184478;
assign addr[16532]= -2106406677;
assign addr[16533]= -2119956737;
assign addr[16534]= -2130817471;
assign addr[16535]= -2138975100;
assign addr[16536]= -2144419275;
assign addr[16537]= -2147143090;
assign addr[16538]= -2147143090;
assign addr[16539]= -2144419275;
assign addr[16540]= -2138975100;
assign addr[16541]= -2130817471;
assign addr[16542]= -2119956737;
assign addr[16543]= -2106406677;
assign addr[16544]= -2090184478;
assign addr[16545]= -2071310720;
assign addr[16546]= -2049809346;
assign addr[16547]= -2025707632;
assign addr[16548]= -1999036154;
assign addr[16549]= -1969828744;
assign addr[16550]= -1938122457;
assign addr[16551]= -1903957513;
assign addr[16552]= -1867377253;
assign addr[16553]= -1828428082;
assign addr[16554]= -1787159411;
assign addr[16555]= -1743623590;
assign addr[16556]= -1697875851;
assign addr[16557]= -1649974225;
assign addr[16558]= -1599979481;
assign addr[16559]= -1547955041;
assign addr[16560]= -1493966902;
assign addr[16561]= -1438083551;
assign addr[16562]= -1380375881;
assign addr[16563]= -1320917099;
assign addr[16564]= -1259782632;
assign addr[16565]= -1197050035;
assign addr[16566]= -1132798888;
assign addr[16567]= -1067110699;
assign addr[16568]= -1000068799;
assign addr[16569]= -931758235;
assign addr[16570]= -862265664;
assign addr[16571]= -791679244;
assign addr[16572]= -720088517;
assign addr[16573]= -647584304;
assign addr[16574]= -574258580;
assign addr[16575]= -500204365;
assign addr[16576]= -425515602;
assign addr[16577]= -350287041;
assign addr[16578]= -274614114;
assign addr[16579]= -198592817;
assign addr[16580]= -122319591;
assign addr[16581]= -45891193;
assign addr[16582]= 30595422;
assign addr[16583]= 107043224;
assign addr[16584]= 183355234;
assign addr[16585]= 259434643;
assign addr[16586]= 335184940;
assign addr[16587]= 410510029;
assign addr[16588]= 485314355;
assign addr[16589]= 559503022;
assign addr[16590]= 632981917;
assign addr[16591]= 705657826;
assign addr[16592]= 777438554;
assign addr[16593]= 848233042;
assign addr[16594]= 917951481;
assign addr[16595]= 986505429;
assign addr[16596]= 1053807919;
assign addr[16597]= 1119773573;
assign addr[16598]= 1184318708;
assign addr[16599]= 1247361445;
assign addr[16600]= 1308821808;
assign addr[16601]= 1368621831;
assign addr[16602]= 1426685652;
assign addr[16603]= 1482939614;
assign addr[16604]= 1537312353;
assign addr[16605]= 1589734894;
assign addr[16606]= 1640140734;
assign addr[16607]= 1688465931;
assign addr[16608]= 1734649179;
assign addr[16609]= 1778631892;
assign addr[16610]= 1820358275;
assign addr[16611]= 1859775393;
assign addr[16612]= 1896833245;
assign addr[16613]= 1931484818;
assign addr[16614]= 1963686155;
assign addr[16615]= 1993396407;
assign addr[16616]= 2020577882;
assign addr[16617]= 2045196100;
assign addr[16618]= 2067219829;
assign addr[16619]= 2086621133;
assign addr[16620]= 2103375398;
assign addr[16621]= 2117461370;
assign addr[16622]= 2128861181;
assign addr[16623]= 2137560369;
assign addr[16624]= 2143547897;
assign addr[16625]= 2146816171;
assign addr[16626]= 2147361045;
assign addr[16627]= 2145181827;
assign addr[16628]= 2140281282;
assign addr[16629]= 2132665626;
assign addr[16630]= 2122344521;
assign addr[16631]= 2109331059;
assign addr[16632]= 2093641749;
assign addr[16633]= 2075296495;
assign addr[16634]= 2054318569;
assign addr[16635]= 2030734582;
assign addr[16636]= 2004574453;
assign addr[16637]= 1975871368;
assign addr[16638]= 1944661739;
assign addr[16639]= 1910985158;
assign addr[16640]= 1874884346;
assign addr[16641]= 1836405100;
assign addr[16642]= 1795596234;
assign addr[16643]= 1752509516;
assign addr[16644]= 1707199606;
assign addr[16645]= 1659723983;
assign addr[16646]= 1610142873;
assign addr[16647]= 1558519173;
assign addr[16648]= 1504918373;
assign addr[16649]= 1449408469;
assign addr[16650]= 1392059879;
assign addr[16651]= 1332945355;
assign addr[16652]= 1272139887;
assign addr[16653]= 1209720613;
assign addr[16654]= 1145766716;
assign addr[16655]= 1080359326;
assign addr[16656]= 1013581418;
assign addr[16657]= 945517704;
assign addr[16658]= 876254528;
assign addr[16659]= 805879757;
assign addr[16660]= 734482665;
assign addr[16661]= 662153826;
assign addr[16662]= 588984994;
assign addr[16663]= 515068990;
assign addr[16664]= 440499581;
assign addr[16665]= 365371365;
assign addr[16666]= 289779648;
assign addr[16667]= 213820322;
assign addr[16668]= 137589750;
assign addr[16669]= 61184634;
assign addr[16670]= -15298099;
assign addr[16671]= -91761426;
assign addr[16672]= -168108346;
assign addr[16673]= -244242007;
assign addr[16674]= -320065829;
assign addr[16675]= -395483624;
assign addr[16676]= -470399716;
assign addr[16677]= -544719071;
assign addr[16678]= -618347408;
assign addr[16679]= -691191324;
assign addr[16680]= -763158411;
assign addr[16681]= -834157373;
assign addr[16682]= -904098143;
assign addr[16683]= -972891995;
assign addr[16684]= -1040451659;
assign addr[16685]= -1106691431;
assign addr[16686]= -1171527280;
assign addr[16687]= -1234876957;
assign addr[16688]= -1296660098;
assign addr[16689]= -1356798326;
assign addr[16690]= -1415215352;
assign addr[16691]= -1471837070;
assign addr[16692]= -1526591649;
assign addr[16693]= -1579409630;
assign addr[16694]= -1630224009;
assign addr[16695]= -1678970324;
assign addr[16696]= -1725586737;
assign addr[16697]= -1770014111;
assign addr[16698]= -1812196087;
assign addr[16699]= -1852079154;
assign addr[16700]= -1889612716;
assign addr[16701]= -1924749160;
assign addr[16702]= -1957443913;
assign addr[16703]= -1987655498;
assign addr[16704]= -2015345591;
assign addr[16705]= -2040479063;
assign addr[16706]= -2063024031;
assign addr[16707]= -2082951896;
assign addr[16708]= -2100237377;
assign addr[16709]= -2114858546;
assign addr[16710]= -2126796855;
assign addr[16711]= -2136037160;
assign addr[16712]= -2142567738;
assign addr[16713]= -2146380306;
assign addr[16714]= -2147470025;
assign addr[16715]= -2145835515;
assign addr[16716]= -2141478848;
assign addr[16717]= -2134405552;
assign addr[16718]= -2124624598;
assign addr[16719]= -2112148396;
assign addr[16720]= -2096992772;
assign addr[16721]= -2079176953;
assign addr[16722]= -2058723538;
assign addr[16723]= -2035658475;
assign addr[16724]= -2010011024;
assign addr[16725]= -1981813720;
assign addr[16726]= -1951102334;
assign addr[16727]= -1917915825;
assign addr[16728]= -1882296293;
assign addr[16729]= -1844288924;
assign addr[16730]= -1803941934;
assign addr[16731]= -1761306505;
assign addr[16732]= -1716436725;
assign addr[16733]= -1669389513;
assign addr[16734]= -1620224553;
assign addr[16735]= -1569004214;
assign addr[16736]= -1515793473;
assign addr[16737]= -1460659832;
assign addr[16738]= -1403673233;
assign addr[16739]= -1344905966;
assign addr[16740]= -1284432584;
assign addr[16741]= -1222329801;
assign addr[16742]= -1158676398;
assign addr[16743]= -1093553126;
assign addr[16744]= -1027042599;
assign addr[16745]= -959229189;
assign addr[16746]= -890198924;
assign addr[16747]= -820039373;
assign addr[16748]= -748839539;
assign addr[16749]= -676689746;
assign addr[16750]= -603681519;
assign addr[16751]= -529907477;
assign addr[16752]= -455461206;
assign addr[16753]= -380437148;
assign addr[16754]= -304930476;
assign addr[16755]= -229036977;
assign addr[16756]= -152852926;
assign addr[16757]= -76474970;
assign addr[16758]= 0;
assign addr[16759]= 76474970;
assign addr[16760]= 152852926;
assign addr[16761]= 229036977;
assign addr[16762]= 304930476;
assign addr[16763]= 380437148;
assign addr[16764]= 455461206;
assign addr[16765]= 529907477;
assign addr[16766]= 603681519;
assign addr[16767]= 676689746;
assign addr[16768]= 748839539;
assign addr[16769]= 820039373;
assign addr[16770]= 890198924;
assign addr[16771]= 959229189;
assign addr[16772]= 1027042599;
assign addr[16773]= 1093553126;
assign addr[16774]= 1158676398;
assign addr[16775]= 1222329801;
assign addr[16776]= 1284432584;
assign addr[16777]= 1344905966;
assign addr[16778]= 1403673233;
assign addr[16779]= 1460659832;
assign addr[16780]= 1515793473;
assign addr[16781]= 1569004214;
assign addr[16782]= 1620224553;
assign addr[16783]= 1669389513;
assign addr[16784]= 1716436725;
assign addr[16785]= 1761306505;
assign addr[16786]= 1803941934;
assign addr[16787]= 1844288924;
assign addr[16788]= 1882296293;
assign addr[16789]= 1917915825;
assign addr[16790]= 1951102334;
assign addr[16791]= 1981813720;
assign addr[16792]= 2010011024;
assign addr[16793]= 2035658475;
assign addr[16794]= 2058723538;
assign addr[16795]= 2079176953;
assign addr[16796]= 2096992772;
assign addr[16797]= 2112148396;
assign addr[16798]= 2124624598;
assign addr[16799]= 2134405552;
assign addr[16800]= 2141478848;
assign addr[16801]= 2145835515;
assign addr[16802]= 2147470025;
assign addr[16803]= 2146380306;
assign addr[16804]= 2142567738;
assign addr[16805]= 2136037160;
assign addr[16806]= 2126796855;
assign addr[16807]= 2114858546;
assign addr[16808]= 2100237377;
assign addr[16809]= 2082951896;
assign addr[16810]= 2063024031;
assign addr[16811]= 2040479063;
assign addr[16812]= 2015345591;
assign addr[16813]= 1987655498;
assign addr[16814]= 1957443913;
assign addr[16815]= 1924749160;
assign addr[16816]= 1889612716;
assign addr[16817]= 1852079154;
assign addr[16818]= 1812196087;
assign addr[16819]= 1770014111;
assign addr[16820]= 1725586737;
assign addr[16821]= 1678970324;
assign addr[16822]= 1630224009;
assign addr[16823]= 1579409630;
assign addr[16824]= 1526591649;
assign addr[16825]= 1471837070;
assign addr[16826]= 1415215352;
assign addr[16827]= 1356798326;
assign addr[16828]= 1296660098;
assign addr[16829]= 1234876957;
assign addr[16830]= 1171527280;
assign addr[16831]= 1106691431;
assign addr[16832]= 1040451659;
assign addr[16833]= 972891995;
assign addr[16834]= 904098143;
assign addr[16835]= 834157373;
assign addr[16836]= 763158411;
assign addr[16837]= 691191324;
assign addr[16838]= 618347408;
assign addr[16839]= 544719071;
assign addr[16840]= 470399716;
assign addr[16841]= 395483624;
assign addr[16842]= 320065829;
assign addr[16843]= 244242007;
assign addr[16844]= 168108346;
assign addr[16845]= 91761426;
assign addr[16846]= 15298099;
assign addr[16847]= -61184634;
assign addr[16848]= -137589750;
assign addr[16849]= -213820322;
assign addr[16850]= -289779648;
assign addr[16851]= -365371365;
assign addr[16852]= -440499581;
assign addr[16853]= -515068990;
assign addr[16854]= -588984994;
assign addr[16855]= -662153826;
assign addr[16856]= -734482665;
assign addr[16857]= -805879757;
assign addr[16858]= -876254528;
assign addr[16859]= -945517704;
assign addr[16860]= -1013581418;
assign addr[16861]= -1080359326;
assign addr[16862]= -1145766716;
assign addr[16863]= -1209720613;
assign addr[16864]= -1272139887;
assign addr[16865]= -1332945355;
assign addr[16866]= -1392059879;
assign addr[16867]= -1449408469;
assign addr[16868]= -1504918373;
assign addr[16869]= -1558519173;
assign addr[16870]= -1610142873;
assign addr[16871]= -1659723983;
assign addr[16872]= -1707199606;
assign addr[16873]= -1752509516;
assign addr[16874]= -1795596234;
assign addr[16875]= -1836405100;
assign addr[16876]= -1874884346;
assign addr[16877]= -1910985158;
assign addr[16878]= -1944661739;
assign addr[16879]= -1975871368;
assign addr[16880]= -2004574453;
assign addr[16881]= -2030734582;
assign addr[16882]= -2054318569;
assign addr[16883]= -2075296495;
assign addr[16884]= -2093641749;
assign addr[16885]= -2109331059;
assign addr[16886]= -2122344521;
assign addr[16887]= -2132665626;
assign addr[16888]= -2140281282;
assign addr[16889]= -2145181827;
assign addr[16890]= -2147361045;
assign addr[16891]= -2146816171;
assign addr[16892]= -2143547897;
assign addr[16893]= -2137560369;
assign addr[16894]= -2128861181;
assign addr[16895]= -2117461370;
assign addr[16896]= -2103375398;
assign addr[16897]= -2086621133;
assign addr[16898]= -2067219829;
assign addr[16899]= -2045196100;
assign addr[16900]= -2020577882;
assign addr[16901]= -1993396407;
assign addr[16902]= -1963686155;
assign addr[16903]= -1931484818;
assign addr[16904]= -1896833245;
assign addr[16905]= -1859775393;
assign addr[16906]= -1820358275;
assign addr[16907]= -1778631892;
assign addr[16908]= -1734649179;
assign addr[16909]= -1688465931;
assign addr[16910]= -1640140734;
assign addr[16911]= -1589734894;
assign addr[16912]= -1537312353;
assign addr[16913]= -1482939614;
assign addr[16914]= -1426685652;
assign addr[16915]= -1368621831;
assign addr[16916]= -1308821808;
assign addr[16917]= -1247361445;
assign addr[16918]= -1184318708;
assign addr[16919]= -1119773573;
assign addr[16920]= -1053807919;
assign addr[16921]= -986505429;
assign addr[16922]= -917951481;
assign addr[16923]= -848233042;
assign addr[16924]= -777438554;
assign addr[16925]= -705657826;
assign addr[16926]= -632981917;
assign addr[16927]= -559503022;
assign addr[16928]= -485314355;
assign addr[16929]= -410510029;
assign addr[16930]= -335184940;
assign addr[16931]= -259434643;
assign addr[16932]= -183355234;
assign addr[16933]= -107043224;
assign addr[16934]= -30595422;
assign addr[16935]= 45891193;
assign addr[16936]= 122319591;
assign addr[16937]= 198592817;
assign addr[16938]= 274614114;
assign addr[16939]= 350287041;
assign addr[16940]= 425515602;
assign addr[16941]= 500204365;
assign addr[16942]= 574258580;
assign addr[16943]= 647584304;
assign addr[16944]= 720088517;
assign addr[16945]= 791679244;
assign addr[16946]= 862265664;
assign addr[16947]= 931758235;
assign addr[16948]= 1000068799;
assign addr[16949]= 1067110699;
assign addr[16950]= 1132798888;
assign addr[16951]= 1197050035;
assign addr[16952]= 1259782632;
assign addr[16953]= 1320917099;
assign addr[16954]= 1380375881;
assign addr[16955]= 1438083551;
assign addr[16956]= 1493966902;
assign addr[16957]= 1547955041;
assign addr[16958]= 1599979481;
assign addr[16959]= 1649974225;
assign addr[16960]= 1697875851;
assign addr[16961]= 1743623590;
assign addr[16962]= 1787159411;
assign addr[16963]= 1828428082;
assign addr[16964]= 1867377253;
assign addr[16965]= 1903957513;
assign addr[16966]= 1938122457;
assign addr[16967]= 1969828744;
assign addr[16968]= 1999036154;
assign addr[16969]= 2025707632;
assign addr[16970]= 2049809346;
assign addr[16971]= 2071310720;
assign addr[16972]= 2090184478;
assign addr[16973]= 2106406677;
assign addr[16974]= 2119956737;
assign addr[16975]= 2130817471;
assign addr[16976]= 2138975100;
assign addr[16977]= 2144419275;
assign addr[16978]= 2147143090;
assign addr[16979]= 2147143090;
assign addr[16980]= 2144419275;
assign addr[16981]= 2138975100;
assign addr[16982]= 2130817471;
assign addr[16983]= 2119956737;
assign addr[16984]= 2106406677;
assign addr[16985]= 2090184478;
assign addr[16986]= 2071310720;
assign addr[16987]= 2049809346;
assign addr[16988]= 2025707632;
assign addr[16989]= 1999036154;
assign addr[16990]= 1969828744;
assign addr[16991]= 1938122457;
assign addr[16992]= 1903957513;
assign addr[16993]= 1867377253;
assign addr[16994]= 1828428082;
assign addr[16995]= 1787159411;
assign addr[16996]= 1743623590;
assign addr[16997]= 1697875851;
assign addr[16998]= 1649974225;
assign addr[16999]= 1599979481;
assign addr[17000]= 1547955041;
assign addr[17001]= 1493966902;
assign addr[17002]= 1438083551;
assign addr[17003]= 1380375881;
assign addr[17004]= 1320917099;
assign addr[17005]= 1259782632;
assign addr[17006]= 1197050035;
assign addr[17007]= 1132798888;
assign addr[17008]= 1067110699;
assign addr[17009]= 1000068799;
assign addr[17010]= 931758235;
assign addr[17011]= 862265664;
assign addr[17012]= 791679244;
assign addr[17013]= 720088517;
assign addr[17014]= 647584304;
assign addr[17015]= 574258580;
assign addr[17016]= 500204365;
assign addr[17017]= 425515602;
assign addr[17018]= 350287041;
assign addr[17019]= 274614114;
assign addr[17020]= 198592817;
assign addr[17021]= 122319591;
assign addr[17022]= 45891193;
assign addr[17023]= -30595422;
assign addr[17024]= -107043224;
assign addr[17025]= -183355234;
assign addr[17026]= -259434643;
assign addr[17027]= -335184940;
assign addr[17028]= -410510029;
assign addr[17029]= -485314355;
assign addr[17030]= -559503022;
assign addr[17031]= -632981917;
assign addr[17032]= -705657826;
assign addr[17033]= -777438554;
assign addr[17034]= -848233042;
assign addr[17035]= -917951481;
assign addr[17036]= -986505429;
assign addr[17037]= -1053807919;
assign addr[17038]= -1119773573;
assign addr[17039]= -1184318708;
assign addr[17040]= -1247361445;
assign addr[17041]= -1308821808;
assign addr[17042]= -1368621831;
assign addr[17043]= -1426685652;
assign addr[17044]= -1482939614;
assign addr[17045]= -1537312353;
assign addr[17046]= -1589734894;
assign addr[17047]= -1640140734;
assign addr[17048]= -1688465931;
assign addr[17049]= -1734649179;
assign addr[17050]= -1778631892;
assign addr[17051]= -1820358275;
assign addr[17052]= -1859775393;
assign addr[17053]= -1896833245;
assign addr[17054]= -1931484818;
assign addr[17055]= -1963686155;
assign addr[17056]= -1993396407;
assign addr[17057]= -2020577882;
assign addr[17058]= -2045196100;
assign addr[17059]= -2067219829;
assign addr[17060]= -2086621133;
assign addr[17061]= -2103375398;
assign addr[17062]= -2117461370;
assign addr[17063]= -2128861181;
assign addr[17064]= -2137560369;
assign addr[17065]= -2143547897;
assign addr[17066]= -2146816171;
assign addr[17067]= -2147361045;
assign addr[17068]= -2145181827;
assign addr[17069]= -2140281282;
assign addr[17070]= -2132665626;
assign addr[17071]= -2122344521;
assign addr[17072]= -2109331059;
assign addr[17073]= -2093641749;
assign addr[17074]= -2075296495;
assign addr[17075]= -2054318569;
assign addr[17076]= -2030734582;
assign addr[17077]= -2004574453;
assign addr[17078]= -1975871368;
assign addr[17079]= -1944661739;
assign addr[17080]= -1910985158;
assign addr[17081]= -1874884346;
assign addr[17082]= -1836405100;
assign addr[17083]= -1795596234;
assign addr[17084]= -1752509516;
assign addr[17085]= -1707199606;
assign addr[17086]= -1659723983;
assign addr[17087]= -1610142873;
assign addr[17088]= -1558519173;
assign addr[17089]= -1504918373;
assign addr[17090]= -1449408469;
assign addr[17091]= -1392059879;
assign addr[17092]= -1332945355;
assign addr[17093]= -1272139887;
assign addr[17094]= -1209720613;
assign addr[17095]= -1145766716;
assign addr[17096]= -1080359326;
assign addr[17097]= -1013581418;
assign addr[17098]= -945517704;
assign addr[17099]= -876254528;
assign addr[17100]= -805879757;
assign addr[17101]= -734482665;
assign addr[17102]= -662153826;
assign addr[17103]= -588984994;
assign addr[17104]= -515068990;
assign addr[17105]= -440499581;
assign addr[17106]= -365371365;
assign addr[17107]= -289779648;
assign addr[17108]= -213820322;
assign addr[17109]= -137589750;
assign addr[17110]= -61184634;
assign addr[17111]= 15298099;
assign addr[17112]= 91761426;
assign addr[17113]= 168108346;
assign addr[17114]= 244242007;
assign addr[17115]= 320065829;
assign addr[17116]= 395483624;
assign addr[17117]= 470399716;
assign addr[17118]= 544719071;
assign addr[17119]= 618347408;
assign addr[17120]= 691191324;
assign addr[17121]= 763158411;
assign addr[17122]= 834157373;
assign addr[17123]= 904098143;
assign addr[17124]= 972891995;
assign addr[17125]= 1040451659;
assign addr[17126]= 1106691431;
assign addr[17127]= 1171527280;
assign addr[17128]= 1234876957;
assign addr[17129]= 1296660098;
assign addr[17130]= 1356798326;
assign addr[17131]= 1415215352;
assign addr[17132]= 1471837070;
assign addr[17133]= 1526591649;
assign addr[17134]= 1579409630;
assign addr[17135]= 1630224009;
assign addr[17136]= 1678970324;
assign addr[17137]= 1725586737;
assign addr[17138]= 1770014111;
assign addr[17139]= 1812196087;
assign addr[17140]= 1852079154;
assign addr[17141]= 1889612716;
assign addr[17142]= 1924749160;
assign addr[17143]= 1957443913;
assign addr[17144]= 1987655498;
assign addr[17145]= 2015345591;
assign addr[17146]= 2040479063;
assign addr[17147]= 2063024031;
assign addr[17148]= 2082951896;
assign addr[17149]= 2100237377;
assign addr[17150]= 2114858546;
assign addr[17151]= 2126796855;
assign addr[17152]= 2136037160;
assign addr[17153]= 2142567738;
assign addr[17154]= 2146380306;
assign addr[17155]= 2147470025;
assign addr[17156]= 2145835515;
assign addr[17157]= 2141478848;
assign addr[17158]= 2134405552;
assign addr[17159]= 2124624598;
assign addr[17160]= 2112148396;
assign addr[17161]= 2096992772;
assign addr[17162]= 2079176953;
assign addr[17163]= 2058723538;
assign addr[17164]= 2035658475;
assign addr[17165]= 2010011024;
assign addr[17166]= 1981813720;
assign addr[17167]= 1951102334;
assign addr[17168]= 1917915825;
assign addr[17169]= 1882296293;
assign addr[17170]= 1844288924;
assign addr[17171]= 1803941934;
assign addr[17172]= 1761306505;
assign addr[17173]= 1716436725;
assign addr[17174]= 1669389513;
assign addr[17175]= 1620224553;
assign addr[17176]= 1569004214;
assign addr[17177]= 1515793473;
assign addr[17178]= 1460659832;
assign addr[17179]= 1403673233;
assign addr[17180]= 1344905966;
assign addr[17181]= 1284432584;
assign addr[17182]= 1222329801;
assign addr[17183]= 1158676398;
assign addr[17184]= 1093553126;
assign addr[17185]= 1027042599;
assign addr[17186]= 959229189;
assign addr[17187]= 890198924;
assign addr[17188]= 820039373;
assign addr[17189]= 748839539;
assign addr[17190]= 676689746;
assign addr[17191]= 603681519;
assign addr[17192]= 529907477;
assign addr[17193]= 455461206;
assign addr[17194]= 380437148;
assign addr[17195]= 304930476;
assign addr[17196]= 229036977;
assign addr[17197]= 152852926;
assign addr[17198]= 76474970;
assign addr[17199]= 0;
assign addr[17200]= -76474970;
assign addr[17201]= -152852926;
assign addr[17202]= -229036977;
assign addr[17203]= -304930476;
assign addr[17204]= -380437148;
assign addr[17205]= -455461206;
assign addr[17206]= -529907477;
assign addr[17207]= -603681519;
assign addr[17208]= -676689746;
assign addr[17209]= -748839539;
assign addr[17210]= -820039373;
assign addr[17211]= -890198924;
assign addr[17212]= -959229189;
assign addr[17213]= -1027042599;
assign addr[17214]= -1093553126;
assign addr[17215]= -1158676398;
assign addr[17216]= -1222329801;
assign addr[17217]= -1284432584;
assign addr[17218]= -1344905966;
assign addr[17219]= -1403673233;
assign addr[17220]= -1460659832;
assign addr[17221]= -1515793473;
assign addr[17222]= -1569004214;
assign addr[17223]= -1620224553;
assign addr[17224]= -1669389513;
assign addr[17225]= -1716436725;
assign addr[17226]= -1761306505;
assign addr[17227]= -1803941934;
assign addr[17228]= -1844288924;
assign addr[17229]= -1882296293;
assign addr[17230]= -1917915825;
assign addr[17231]= -1951102334;
assign addr[17232]= -1981813720;
assign addr[17233]= -2010011024;
assign addr[17234]= -2035658475;
assign addr[17235]= -2058723538;
assign addr[17236]= -2079176953;
assign addr[17237]= -2096992772;
assign addr[17238]= -2112148396;
assign addr[17239]= -2124624598;
assign addr[17240]= -2134405552;
assign addr[17241]= -2141478848;
assign addr[17242]= -2145835515;
assign addr[17243]= -2147470025;
assign addr[17244]= -2146380306;
assign addr[17245]= -2142567738;
assign addr[17246]= -2136037160;
assign addr[17247]= -2126796855;
assign addr[17248]= -2114858546;
assign addr[17249]= -2100237377;
assign addr[17250]= -2082951896;
assign addr[17251]= -2063024031;
assign addr[17252]= -2040479063;
assign addr[17253]= -2015345591;
assign addr[17254]= -1987655498;
assign addr[17255]= -1957443913;
assign addr[17256]= -1924749160;
assign addr[17257]= -1889612716;
assign addr[17258]= -1852079154;
assign addr[17259]= -1812196087;
assign addr[17260]= -1770014111;
assign addr[17261]= -1725586737;
assign addr[17262]= -1678970324;
assign addr[17263]= -1630224009;
assign addr[17264]= -1579409630;
assign addr[17265]= -1526591649;
assign addr[17266]= -1471837070;
assign addr[17267]= -1415215352;
assign addr[17268]= -1356798326;
assign addr[17269]= -1296660098;
assign addr[17270]= -1234876957;
assign addr[17271]= -1171527280;
assign addr[17272]= -1106691431;
assign addr[17273]= -1040451659;
assign addr[17274]= -972891995;
assign addr[17275]= -904098143;
assign addr[17276]= -834157373;
assign addr[17277]= -763158411;
assign addr[17278]= -691191324;
assign addr[17279]= -618347408;
assign addr[17280]= -544719071;
assign addr[17281]= -470399716;
assign addr[17282]= -395483624;
assign addr[17283]= -320065829;
assign addr[17284]= -244242007;
assign addr[17285]= -168108346;
assign addr[17286]= -91761426;
assign addr[17287]= -15298099;
assign addr[17288]= 61184634;
assign addr[17289]= 137589750;
assign addr[17290]= 213820322;
assign addr[17291]= 289779648;
assign addr[17292]= 365371365;
assign addr[17293]= 440499581;
assign addr[17294]= 515068990;
assign addr[17295]= 588984994;
assign addr[17296]= 662153826;
assign addr[17297]= 734482665;
assign addr[17298]= 805879757;
assign addr[17299]= 876254528;
assign addr[17300]= 945517704;
assign addr[17301]= 1013581418;
assign addr[17302]= 1080359326;
assign addr[17303]= 1145766716;
assign addr[17304]= 1209720613;
assign addr[17305]= 1272139887;
assign addr[17306]= 1332945355;
assign addr[17307]= 1392059879;
assign addr[17308]= 1449408469;
assign addr[17309]= 1504918373;
assign addr[17310]= 1558519173;
assign addr[17311]= 1610142873;
assign addr[17312]= 1659723983;
assign addr[17313]= 1707199606;
assign addr[17314]= 1752509516;
assign addr[17315]= 1795596234;
assign addr[17316]= 1836405100;
assign addr[17317]= 1874884346;
assign addr[17318]= 1910985158;
assign addr[17319]= 1944661739;
assign addr[17320]= 1975871368;
assign addr[17321]= 2004574453;
assign addr[17322]= 2030734582;
assign addr[17323]= 2054318569;
assign addr[17324]= 2075296495;
assign addr[17325]= 2093641749;
assign addr[17326]= 2109331059;
assign addr[17327]= 2122344521;
assign addr[17328]= 2132665626;
assign addr[17329]= 2140281282;
assign addr[17330]= 2145181827;
assign addr[17331]= 2147361045;
assign addr[17332]= 2146816171;
assign addr[17333]= 2143547897;
assign addr[17334]= 2137560369;
assign addr[17335]= 2128861181;
assign addr[17336]= 2117461370;
assign addr[17337]= 2103375398;
assign addr[17338]= 2086621133;
assign addr[17339]= 2067219829;
assign addr[17340]= 2045196100;
assign addr[17341]= 2020577882;
assign addr[17342]= 1993396407;
assign addr[17343]= 1963686155;
assign addr[17344]= 1931484818;
assign addr[17345]= 1896833245;
assign addr[17346]= 1859775393;
assign addr[17347]= 1820358275;
assign addr[17348]= 1778631892;
assign addr[17349]= 1734649179;
assign addr[17350]= 1688465931;
assign addr[17351]= 1640140734;
assign addr[17352]= 1589734894;
assign addr[17353]= 1537312353;
assign addr[17354]= 1482939614;
assign addr[17355]= 1426685652;
assign addr[17356]= 1368621831;
assign addr[17357]= 1308821808;
assign addr[17358]= 1247361445;
assign addr[17359]= 1184318708;
assign addr[17360]= 1119773573;
assign addr[17361]= 1053807919;
assign addr[17362]= 986505429;
assign addr[17363]= 917951481;
assign addr[17364]= 848233042;
assign addr[17365]= 777438554;
assign addr[17366]= 705657826;
assign addr[17367]= 632981917;
assign addr[17368]= 559503022;
assign addr[17369]= 485314355;
assign addr[17370]= 410510029;
assign addr[17371]= 335184940;
assign addr[17372]= 259434643;
assign addr[17373]= 183355234;
assign addr[17374]= 107043224;
assign addr[17375]= 30595422;
assign addr[17376]= -45891193;
assign addr[17377]= -122319591;
assign addr[17378]= -198592817;
assign addr[17379]= -274614114;
assign addr[17380]= -350287041;
assign addr[17381]= -425515602;
assign addr[17382]= -500204365;
assign addr[17383]= -574258580;
assign addr[17384]= -647584304;
assign addr[17385]= -720088517;
assign addr[17386]= -791679244;
assign addr[17387]= -862265664;
assign addr[17388]= -931758235;
assign addr[17389]= -1000068799;
assign addr[17390]= -1067110699;
assign addr[17391]= -1132798888;
assign addr[17392]= -1197050035;
assign addr[17393]= -1259782632;
assign addr[17394]= -1320917099;
assign addr[17395]= -1380375881;
assign addr[17396]= -1438083551;
assign addr[17397]= -1493966902;
assign addr[17398]= -1547955041;
assign addr[17399]= -1599979481;
assign addr[17400]= -1649974225;
assign addr[17401]= -1697875851;
assign addr[17402]= -1743623590;
assign addr[17403]= -1787159411;
assign addr[17404]= -1828428082;
assign addr[17405]= -1867377253;
assign addr[17406]= -1903957513;
assign addr[17407]= -1938122457;
assign addr[17408]= -1969828744;
assign addr[17409]= -1999036154;
assign addr[17410]= -2025707632;
assign addr[17411]= -2049809346;
assign addr[17412]= -2071310720;
assign addr[17413]= -2090184478;
assign addr[17414]= -2106406677;
assign addr[17415]= -2119956737;
assign addr[17416]= -2130817471;
assign addr[17417]= -2138975100;
assign addr[17418]= -2144419275;
assign addr[17419]= -2147143090;
assign addr[17420]= -2147143090;
assign addr[17421]= -2144419275;
assign addr[17422]= -2138975100;
assign addr[17423]= -2130817471;
assign addr[17424]= -2119956737;
assign addr[17425]= -2106406677;
assign addr[17426]= -2090184478;
assign addr[17427]= -2071310720;
assign addr[17428]= -2049809346;
assign addr[17429]= -2025707632;
assign addr[17430]= -1999036154;
assign addr[17431]= -1969828744;
assign addr[17432]= -1938122457;
assign addr[17433]= -1903957513;
assign addr[17434]= -1867377253;
assign addr[17435]= -1828428082;
assign addr[17436]= -1787159411;
assign addr[17437]= -1743623590;
assign addr[17438]= -1697875851;
assign addr[17439]= -1649974225;
assign addr[17440]= -1599979481;
assign addr[17441]= -1547955041;
assign addr[17442]= -1493966902;
assign addr[17443]= -1438083551;
assign addr[17444]= -1380375881;
assign addr[17445]= -1320917099;
assign addr[17446]= -1259782632;
assign addr[17447]= -1197050035;
assign addr[17448]= -1132798888;
assign addr[17449]= -1067110699;
assign addr[17450]= -1000068799;
assign addr[17451]= -931758235;
assign addr[17452]= -862265664;
assign addr[17453]= -791679244;
assign addr[17454]= -720088517;
assign addr[17455]= -647584304;
assign addr[17456]= -574258580;
assign addr[17457]= -500204365;
assign addr[17458]= -425515602;
assign addr[17459]= -350287041;
assign addr[17460]= -274614114;
assign addr[17461]= -198592817;
assign addr[17462]= -122319591;
assign addr[17463]= -45891193;
assign addr[17464]= 30595422;
assign addr[17465]= 107043224;
assign addr[17466]= 183355234;
assign addr[17467]= 259434643;
assign addr[17468]= 335184940;
assign addr[17469]= 410510029;
assign addr[17470]= 485314355;
assign addr[17471]= 559503022;
assign addr[17472]= 632981917;
assign addr[17473]= 705657826;
assign addr[17474]= 777438554;
assign addr[17475]= 848233042;
assign addr[17476]= 917951481;
assign addr[17477]= 986505429;
assign addr[17478]= 1053807919;
assign addr[17479]= 1119773573;
assign addr[17480]= 1184318708;
assign addr[17481]= 1247361445;
assign addr[17482]= 1308821808;
assign addr[17483]= 1368621831;
assign addr[17484]= 1426685652;
assign addr[17485]= 1482939614;
assign addr[17486]= 1537312353;
assign addr[17487]= 1589734894;
assign addr[17488]= 1640140734;
assign addr[17489]= 1688465931;
assign addr[17490]= 1734649179;
assign addr[17491]= 1778631892;
assign addr[17492]= 1820358275;
assign addr[17493]= 1859775393;
assign addr[17494]= 1896833245;
assign addr[17495]= 1931484818;
assign addr[17496]= 1963686155;
assign addr[17497]= 1993396407;
assign addr[17498]= 2020577882;
assign addr[17499]= 2045196100;
assign addr[17500]= 2067219829;
assign addr[17501]= 2086621133;
assign addr[17502]= 2103375398;
assign addr[17503]= 2117461370;
assign addr[17504]= 2128861181;
assign addr[17505]= 2137560369;
assign addr[17506]= 2143547897;
assign addr[17507]= 2146816171;
assign addr[17508]= 2147361045;
assign addr[17509]= 2145181827;
assign addr[17510]= 2140281282;
assign addr[17511]= 2132665626;
assign addr[17512]= 2122344521;
assign addr[17513]= 2109331059;
assign addr[17514]= 2093641749;
assign addr[17515]= 2075296495;
assign addr[17516]= 2054318569;
assign addr[17517]= 2030734582;
assign addr[17518]= 2004574453;
assign addr[17519]= 1975871368;
assign addr[17520]= 1944661739;
assign addr[17521]= 1910985158;
assign addr[17522]= 1874884346;
assign addr[17523]= 1836405100;
assign addr[17524]= 1795596234;
assign addr[17525]= 1752509516;
assign addr[17526]= 1707199606;
assign addr[17527]= 1659723983;
assign addr[17528]= 1610142873;
assign addr[17529]= 1558519173;
assign addr[17530]= 1504918373;
assign addr[17531]= 1449408469;
assign addr[17532]= 1392059879;
assign addr[17533]= 1332945355;
assign addr[17534]= 1272139887;
assign addr[17535]= 1209720613;
assign addr[17536]= 1145766716;
assign addr[17537]= 1080359326;
assign addr[17538]= 1013581418;
assign addr[17539]= 945517704;
assign addr[17540]= 876254528;
assign addr[17541]= 805879757;
assign addr[17542]= 734482665;
assign addr[17543]= 662153826;
assign addr[17544]= 588984994;
assign addr[17545]= 515068990;
assign addr[17546]= 440499581;
assign addr[17547]= 365371365;
assign addr[17548]= 289779648;
assign addr[17549]= 213820322;
assign addr[17550]= 137589750;
assign addr[17551]= 61184634;
assign addr[17552]= -15298099;
assign addr[17553]= -91761426;
assign addr[17554]= -168108346;
assign addr[17555]= -244242007;
assign addr[17556]= -320065829;
assign addr[17557]= -395483624;
assign addr[17558]= -470399716;
assign addr[17559]= -544719071;
assign addr[17560]= -618347408;
assign addr[17561]= -691191324;
assign addr[17562]= -763158411;
assign addr[17563]= -834157373;
assign addr[17564]= -904098143;
assign addr[17565]= -972891995;
assign addr[17566]= -1040451659;
assign addr[17567]= -1106691431;
assign addr[17568]= -1171527280;
assign addr[17569]= -1234876957;
assign addr[17570]= -1296660098;
assign addr[17571]= -1356798326;
assign addr[17572]= -1415215352;
assign addr[17573]= -1471837070;
assign addr[17574]= -1526591649;
assign addr[17575]= -1579409630;
assign addr[17576]= -1630224009;
assign addr[17577]= -1678970324;
assign addr[17578]= -1725586737;
assign addr[17579]= -1770014111;
assign addr[17580]= -1812196087;
assign addr[17581]= -1852079154;
assign addr[17582]= -1889612716;
assign addr[17583]= -1924749160;
assign addr[17584]= -1957443913;
assign addr[17585]= -1987655498;
assign addr[17586]= -2015345591;
assign addr[17587]= -2040479063;
assign addr[17588]= -2063024031;
assign addr[17589]= -2082951896;
assign addr[17590]= -2100237377;
assign addr[17591]= -2114858546;
assign addr[17592]= -2126796855;
assign addr[17593]= -2136037160;
assign addr[17594]= -2142567738;
assign addr[17595]= -2146380306;
assign addr[17596]= -2147470025;
assign addr[17597]= -2145835515;
assign addr[17598]= -2141478848;
assign addr[17599]= -2134405552;
assign addr[17600]= -2124624598;
assign addr[17601]= -2112148396;
assign addr[17602]= -2096992772;
assign addr[17603]= -2079176953;
assign addr[17604]= -2058723538;
assign addr[17605]= -2035658475;
assign addr[17606]= -2010011024;
assign addr[17607]= -1981813720;
assign addr[17608]= -1951102334;
assign addr[17609]= -1917915825;
assign addr[17610]= -1882296293;
assign addr[17611]= -1844288924;
assign addr[17612]= -1803941934;
assign addr[17613]= -1761306505;
assign addr[17614]= -1716436725;
assign addr[17615]= -1669389513;
assign addr[17616]= -1620224553;
assign addr[17617]= -1569004214;
assign addr[17618]= -1515793473;
assign addr[17619]= -1460659832;
assign addr[17620]= -1403673233;
assign addr[17621]= -1344905966;
assign addr[17622]= -1284432584;
assign addr[17623]= -1222329801;
assign addr[17624]= -1158676398;
assign addr[17625]= -1093553126;
assign addr[17626]= -1027042599;
assign addr[17627]= -959229189;
assign addr[17628]= -890198924;
assign addr[17629]= -820039373;
assign addr[17630]= -748839539;
assign addr[17631]= -676689746;
assign addr[17632]= -603681519;
assign addr[17633]= -529907477;
assign addr[17634]= -455461206;
assign addr[17635]= -380437148;
assign addr[17636]= -304930476;
assign addr[17637]= -229036977;
assign addr[17638]= -152852926;
assign addr[17639]= -76474970;
assign addr[17640]= 0;
assign addr[17641]= 76474970;
assign addr[17642]= 152852926;
assign addr[17643]= 229036977;
assign addr[17644]= 304930476;
assign addr[17645]= 380437148;
assign addr[17646]= 455461206;
assign addr[17647]= 529907477;
assign addr[17648]= 603681519;
assign addr[17649]= 676689746;
assign addr[17650]= 748839539;
assign addr[17651]= 820039373;
assign addr[17652]= 890198924;
assign addr[17653]= 959229189;
assign addr[17654]= 1027042599;
assign addr[17655]= 1093553126;
assign addr[17656]= 1158676398;
assign addr[17657]= 1222329801;
assign addr[17658]= 1284432584;
assign addr[17659]= 1344905966;
assign addr[17660]= 1403673233;
assign addr[17661]= 1460659832;
assign addr[17662]= 1515793473;
assign addr[17663]= 1569004214;
assign addr[17664]= 1620224553;
assign addr[17665]= 1669389513;
assign addr[17666]= 1716436725;
assign addr[17667]= 1761306505;
assign addr[17668]= 1803941934;
assign addr[17669]= 1844288924;
assign addr[17670]= 1882296293;
assign addr[17671]= 1917915825;
assign addr[17672]= 1951102334;
assign addr[17673]= 1981813720;
assign addr[17674]= 2010011024;
assign addr[17675]= 2035658475;
assign addr[17676]= 2058723538;
assign addr[17677]= 2079176953;
assign addr[17678]= 2096992772;
assign addr[17679]= 2112148396;
assign addr[17680]= 2124624598;
assign addr[17681]= 2134405552;
assign addr[17682]= 2141478848;
assign addr[17683]= 2145835515;
assign addr[17684]= 2147470025;
assign addr[17685]= 2146380306;
assign addr[17686]= 2142567738;
assign addr[17687]= 2136037160;
assign addr[17688]= 2126796855;
assign addr[17689]= 2114858546;
assign addr[17690]= 2100237377;
assign addr[17691]= 2082951896;
assign addr[17692]= 2063024031;
assign addr[17693]= 2040479063;
assign addr[17694]= 2015345591;
assign addr[17695]= 1987655498;
assign addr[17696]= 1957443913;
assign addr[17697]= 1924749160;
assign addr[17698]= 1889612716;
assign addr[17699]= 1852079154;
assign addr[17700]= 1812196087;
assign addr[17701]= 1770014111;
assign addr[17702]= 1725586737;
assign addr[17703]= 1678970324;
assign addr[17704]= 1630224009;
assign addr[17705]= 1579409630;
assign addr[17706]= 1526591649;
assign addr[17707]= 1471837070;
assign addr[17708]= 1415215352;
assign addr[17709]= 1356798326;
assign addr[17710]= 1296660098;
assign addr[17711]= 1234876957;
assign addr[17712]= 1171527280;
assign addr[17713]= 1106691431;
assign addr[17714]= 1040451659;
assign addr[17715]= 972891995;
assign addr[17716]= 904098143;
assign addr[17717]= 834157373;
assign addr[17718]= 763158411;
assign addr[17719]= 691191324;
assign addr[17720]= 618347408;
assign addr[17721]= 544719071;
assign addr[17722]= 470399716;
assign addr[17723]= 395483624;
assign addr[17724]= 320065829;
assign addr[17725]= 244242007;
assign addr[17726]= 168108346;
assign addr[17727]= 91761426;
assign addr[17728]= 15298099;
assign addr[17729]= -61184634;
assign addr[17730]= -137589750;
assign addr[17731]= -213820322;
assign addr[17732]= -289779648;
assign addr[17733]= -365371365;
assign addr[17734]= -440499581;
assign addr[17735]= -515068990;
assign addr[17736]= -588984994;
assign addr[17737]= -662153826;
assign addr[17738]= -734482665;
assign addr[17739]= -805879757;
assign addr[17740]= -876254528;
assign addr[17741]= -945517704;
assign addr[17742]= -1013581418;
assign addr[17743]= -1080359326;
assign addr[17744]= -1145766716;
assign addr[17745]= -1209720613;
assign addr[17746]= -1272139887;
assign addr[17747]= -1332945355;
assign addr[17748]= -1392059879;
assign addr[17749]= -1449408469;
assign addr[17750]= -1504918373;
assign addr[17751]= -1558519173;
assign addr[17752]= -1610142873;
assign addr[17753]= -1659723983;
assign addr[17754]= -1707199606;
assign addr[17755]= -1752509516;
assign addr[17756]= -1795596234;
assign addr[17757]= -1836405100;
assign addr[17758]= -1874884346;
assign addr[17759]= -1910985158;
assign addr[17760]= -1944661739;
assign addr[17761]= -1975871368;
assign addr[17762]= -2004574453;
assign addr[17763]= -2030734582;
assign addr[17764]= -2054318569;
assign addr[17765]= -2075296495;
assign addr[17766]= -2093641749;
assign addr[17767]= -2109331059;
assign addr[17768]= -2122344521;
assign addr[17769]= -2132665626;
assign addr[17770]= -2140281282;
assign addr[17771]= -2145181827;
assign addr[17772]= -2147361045;
assign addr[17773]= -2146816171;
assign addr[17774]= -2143547897;
assign addr[17775]= -2137560369;
assign addr[17776]= -2128861181;
assign addr[17777]= -2117461370;
assign addr[17778]= -2103375398;
assign addr[17779]= -2086621133;
assign addr[17780]= -2067219829;
assign addr[17781]= -2045196100;
assign addr[17782]= -2020577882;
assign addr[17783]= -1993396407;
assign addr[17784]= -1963686155;
assign addr[17785]= -1931484818;
assign addr[17786]= -1896833245;
assign addr[17787]= -1859775393;
assign addr[17788]= -1820358275;
assign addr[17789]= -1778631892;
assign addr[17790]= -1734649179;
assign addr[17791]= -1688465931;
assign addr[17792]= -1640140734;
assign addr[17793]= -1589734894;
assign addr[17794]= -1537312353;
assign addr[17795]= -1482939614;
assign addr[17796]= -1426685652;
assign addr[17797]= -1368621831;
assign addr[17798]= -1308821808;
assign addr[17799]= -1247361445;
assign addr[17800]= -1184318708;
assign addr[17801]= -1119773573;
assign addr[17802]= -1053807919;
assign addr[17803]= -986505429;
assign addr[17804]= -917951481;
assign addr[17805]= -848233042;
assign addr[17806]= -777438554;
assign addr[17807]= -705657826;
assign addr[17808]= -632981917;
assign addr[17809]= -559503022;
assign addr[17810]= -485314355;
assign addr[17811]= -410510029;
assign addr[17812]= -335184940;
assign addr[17813]= -259434643;
assign addr[17814]= -183355234;
assign addr[17815]= -107043224;
assign addr[17816]= -30595422;
assign addr[17817]= 45891193;
assign addr[17818]= 122319591;
assign addr[17819]= 198592817;
assign addr[17820]= 274614114;
assign addr[17821]= 350287041;
assign addr[17822]= 425515602;
assign addr[17823]= 500204365;
assign addr[17824]= 574258580;
assign addr[17825]= 647584304;
assign addr[17826]= 720088517;
assign addr[17827]= 791679244;
assign addr[17828]= 862265664;
assign addr[17829]= 931758235;
assign addr[17830]= 1000068799;
assign addr[17831]= 1067110699;
assign addr[17832]= 1132798888;
assign addr[17833]= 1197050035;
assign addr[17834]= 1259782632;
assign addr[17835]= 1320917099;
assign addr[17836]= 1380375881;
assign addr[17837]= 1438083551;
assign addr[17838]= 1493966902;
assign addr[17839]= 1547955041;
assign addr[17840]= 1599979481;
assign addr[17841]= 1649974225;
assign addr[17842]= 1697875851;
assign addr[17843]= 1743623590;
assign addr[17844]= 1787159411;
assign addr[17845]= 1828428082;
assign addr[17846]= 1867377253;
assign addr[17847]= 1903957513;
assign addr[17848]= 1938122457;
assign addr[17849]= 1969828744;
assign addr[17850]= 1999036154;
assign addr[17851]= 2025707632;
assign addr[17852]= 2049809346;
assign addr[17853]= 2071310720;
assign addr[17854]= 2090184478;
assign addr[17855]= 2106406677;
assign addr[17856]= 2119956737;
assign addr[17857]= 2130817471;
assign addr[17858]= 2138975100;
assign addr[17859]= 2144419275;
assign addr[17860]= 2147143090;
assign addr[17861]= 2147143090;
assign addr[17862]= 2144419275;
assign addr[17863]= 2138975100;
assign addr[17864]= 2130817471;
assign addr[17865]= 2119956737;
assign addr[17866]= 2106406677;
assign addr[17867]= 2090184478;
assign addr[17868]= 2071310720;
assign addr[17869]= 2049809346;
assign addr[17870]= 2025707632;
assign addr[17871]= 1999036154;
assign addr[17872]= 1969828744;
assign addr[17873]= 1938122457;
assign addr[17874]= 1903957513;
assign addr[17875]= 1867377253;
assign addr[17876]= 1828428082;
assign addr[17877]= 1787159411;
assign addr[17878]= 1743623590;
assign addr[17879]= 1697875851;
assign addr[17880]= 1649974225;
assign addr[17881]= 1599979481;
assign addr[17882]= 1547955041;
assign addr[17883]= 1493966902;
assign addr[17884]= 1438083551;
assign addr[17885]= 1380375881;
assign addr[17886]= 1320917099;
assign addr[17887]= 1259782632;
assign addr[17888]= 1197050035;
assign addr[17889]= 1132798888;
assign addr[17890]= 1067110699;
assign addr[17891]= 1000068799;
assign addr[17892]= 931758235;
assign addr[17893]= 862265664;
assign addr[17894]= 791679244;
assign addr[17895]= 720088517;
assign addr[17896]= 647584304;
assign addr[17897]= 574258580;
assign addr[17898]= 500204365;
assign addr[17899]= 425515602;
assign addr[17900]= 350287041;
assign addr[17901]= 274614114;
assign addr[17902]= 198592817;
assign addr[17903]= 122319591;
assign addr[17904]= 45891193;
assign addr[17905]= -30595422;
assign addr[17906]= -107043224;
assign addr[17907]= -183355234;
assign addr[17908]= -259434643;
assign addr[17909]= -335184940;
assign addr[17910]= -410510029;
assign addr[17911]= -485314355;
assign addr[17912]= -559503022;
assign addr[17913]= -632981917;
assign addr[17914]= -705657826;
assign addr[17915]= -777438554;
assign addr[17916]= -848233042;
assign addr[17917]= -917951481;
assign addr[17918]= -986505429;
assign addr[17919]= -1053807919;
assign addr[17920]= -1119773573;
assign addr[17921]= -1184318708;
assign addr[17922]= -1247361445;
assign addr[17923]= -1308821808;
assign addr[17924]= -1368621831;
assign addr[17925]= -1426685652;
assign addr[17926]= -1482939614;
assign addr[17927]= -1537312353;
assign addr[17928]= -1589734894;
assign addr[17929]= -1640140734;
assign addr[17930]= -1688465931;
assign addr[17931]= -1734649179;
assign addr[17932]= -1778631892;
assign addr[17933]= -1820358275;
assign addr[17934]= -1859775393;
assign addr[17935]= -1896833245;
assign addr[17936]= -1931484818;
assign addr[17937]= -1963686155;
assign addr[17938]= -1993396407;
assign addr[17939]= -2020577882;
assign addr[17940]= -2045196100;
assign addr[17941]= -2067219829;
assign addr[17942]= -2086621133;
assign addr[17943]= -2103375398;
assign addr[17944]= -2117461370;
assign addr[17945]= -2128861181;
assign addr[17946]= -2137560369;
assign addr[17947]= -2143547897;
assign addr[17948]= -2146816171;
assign addr[17949]= -2147361045;
assign addr[17950]= -2145181827;
assign addr[17951]= -2140281282;
assign addr[17952]= -2132665626;
assign addr[17953]= -2122344521;
assign addr[17954]= -2109331059;
assign addr[17955]= -2093641749;
assign addr[17956]= -2075296495;
assign addr[17957]= -2054318569;
assign addr[17958]= -2030734582;
assign addr[17959]= -2004574453;
assign addr[17960]= -1975871368;
assign addr[17961]= -1944661739;
assign addr[17962]= -1910985158;
assign addr[17963]= -1874884346;
assign addr[17964]= -1836405100;
assign addr[17965]= -1795596234;
assign addr[17966]= -1752509516;
assign addr[17967]= -1707199606;
assign addr[17968]= -1659723983;
assign addr[17969]= -1610142873;
assign addr[17970]= -1558519173;
assign addr[17971]= -1504918373;
assign addr[17972]= -1449408469;
assign addr[17973]= -1392059879;
assign addr[17974]= -1332945355;
assign addr[17975]= -1272139887;
assign addr[17976]= -1209720613;
assign addr[17977]= -1145766716;
assign addr[17978]= -1080359326;
assign addr[17979]= -1013581418;
assign addr[17980]= -945517704;
assign addr[17981]= -876254528;
assign addr[17982]= -805879757;
assign addr[17983]= -734482665;
assign addr[17984]= -662153826;
assign addr[17985]= -588984994;
assign addr[17986]= -515068990;
assign addr[17987]= -440499581;
assign addr[17988]= -365371365;
assign addr[17989]= -289779648;
assign addr[17990]= -213820322;
assign addr[17991]= -137589750;
assign addr[17992]= -61184634;
assign addr[17993]= 15298099;
assign addr[17994]= 91761426;
assign addr[17995]= 168108346;
assign addr[17996]= 244242007;
assign addr[17997]= 320065829;
assign addr[17998]= 395483624;
assign addr[17999]= 470399716;
assign addr[18000]= 544719071;
assign addr[18001]= 618347408;
assign addr[18002]= 691191324;
assign addr[18003]= 763158411;
assign addr[18004]= 834157373;
assign addr[18005]= 904098143;
assign addr[18006]= 972891995;
assign addr[18007]= 1040451659;
assign addr[18008]= 1106691431;
assign addr[18009]= 1171527280;
assign addr[18010]= 1234876957;
assign addr[18011]= 1296660098;
assign addr[18012]= 1356798326;
assign addr[18013]= 1415215352;
assign addr[18014]= 1471837070;
assign addr[18015]= 1526591649;
assign addr[18016]= 1579409630;
assign addr[18017]= 1630224009;
assign addr[18018]= 1678970324;
assign addr[18019]= 1725586737;
assign addr[18020]= 1770014111;
assign addr[18021]= 1812196087;
assign addr[18022]= 1852079154;
assign addr[18023]= 1889612716;
assign addr[18024]= 1924749160;
assign addr[18025]= 1957443913;
assign addr[18026]= 1987655498;
assign addr[18027]= 2015345591;
assign addr[18028]= 2040479063;
assign addr[18029]= 2063024031;
assign addr[18030]= 2082951896;
assign addr[18031]= 2100237377;
assign addr[18032]= 2114858546;
assign addr[18033]= 2126796855;
assign addr[18034]= 2136037160;
assign addr[18035]= 2142567738;
assign addr[18036]= 2146380306;
assign addr[18037]= 2147470025;
assign addr[18038]= 2145835515;
assign addr[18039]= 2141478848;
assign addr[18040]= 2134405552;
assign addr[18041]= 2124624598;
assign addr[18042]= 2112148396;
assign addr[18043]= 2096992772;
assign addr[18044]= 2079176953;
assign addr[18045]= 2058723538;
assign addr[18046]= 2035658475;
assign addr[18047]= 2010011024;
assign addr[18048]= 1981813720;
assign addr[18049]= 1951102334;
assign addr[18050]= 1917915825;
assign addr[18051]= 1882296293;
assign addr[18052]= 1844288924;
assign addr[18053]= 1803941934;
assign addr[18054]= 1761306505;
assign addr[18055]= 1716436725;
assign addr[18056]= 1669389513;
assign addr[18057]= 1620224553;
assign addr[18058]= 1569004214;
assign addr[18059]= 1515793473;
assign addr[18060]= 1460659832;
assign addr[18061]= 1403673233;
assign addr[18062]= 1344905966;
assign addr[18063]= 1284432584;
assign addr[18064]= 1222329801;
assign addr[18065]= 1158676398;
assign addr[18066]= 1093553126;
assign addr[18067]= 1027042599;
assign addr[18068]= 959229189;
assign addr[18069]= 890198924;
assign addr[18070]= 820039373;
assign addr[18071]= 748839539;
assign addr[18072]= 676689746;
assign addr[18073]= 603681519;
assign addr[18074]= 529907477;
assign addr[18075]= 455461206;
assign addr[18076]= 380437148;
assign addr[18077]= 304930476;
assign addr[18078]= 229036977;
assign addr[18079]= 152852926;
assign addr[18080]= 76474970;
assign addr[18081]= 0;
assign addr[18082]= -76474970;
assign addr[18083]= -152852926;
assign addr[18084]= -229036977;
assign addr[18085]= -304930476;
assign addr[18086]= -380437148;
assign addr[18087]= -455461206;
assign addr[18088]= -529907477;
assign addr[18089]= -603681519;
assign addr[18090]= -676689746;
assign addr[18091]= -748839539;
assign addr[18092]= -820039373;
assign addr[18093]= -890198924;
assign addr[18094]= -959229189;
assign addr[18095]= -1027042599;
assign addr[18096]= -1093553126;
assign addr[18097]= -1158676398;
assign addr[18098]= -1222329801;
assign addr[18099]= -1284432584;
assign addr[18100]= -1344905966;
assign addr[18101]= -1403673233;
assign addr[18102]= -1460659832;
assign addr[18103]= -1515793473;
assign addr[18104]= -1569004214;
assign addr[18105]= -1620224553;
assign addr[18106]= -1669389513;
assign addr[18107]= -1716436725;
assign addr[18108]= -1761306505;
assign addr[18109]= -1803941934;
assign addr[18110]= -1844288924;
assign addr[18111]= -1882296293;
assign addr[18112]= -1917915825;
assign addr[18113]= -1951102334;
assign addr[18114]= -1981813720;
assign addr[18115]= -2010011024;
assign addr[18116]= -2035658475;
assign addr[18117]= -2058723538;
assign addr[18118]= -2079176953;
assign addr[18119]= -2096992772;
assign addr[18120]= -2112148396;
assign addr[18121]= -2124624598;
assign addr[18122]= -2134405552;
assign addr[18123]= -2141478848;
assign addr[18124]= -2145835515;
assign addr[18125]= -2147470025;
assign addr[18126]= -2146380306;
assign addr[18127]= -2142567738;
assign addr[18128]= -2136037160;
assign addr[18129]= -2126796855;
assign addr[18130]= -2114858546;
assign addr[18131]= -2100237377;
assign addr[18132]= -2082951896;
assign addr[18133]= -2063024031;
assign addr[18134]= -2040479063;
assign addr[18135]= -2015345591;
assign addr[18136]= -1987655498;
assign addr[18137]= -1957443913;
assign addr[18138]= -1924749160;
assign addr[18139]= -1889612716;
assign addr[18140]= -1852079154;
assign addr[18141]= -1812196087;
assign addr[18142]= -1770014111;
assign addr[18143]= -1725586737;
assign addr[18144]= -1678970324;
assign addr[18145]= -1630224009;
assign addr[18146]= -1579409630;
assign addr[18147]= -1526591649;
assign addr[18148]= -1471837070;
assign addr[18149]= -1415215352;
assign addr[18150]= -1356798326;
assign addr[18151]= -1296660098;
assign addr[18152]= -1234876957;
assign addr[18153]= -1171527280;
assign addr[18154]= -1106691431;
assign addr[18155]= -1040451659;
assign addr[18156]= -972891995;
assign addr[18157]= -904098143;
assign addr[18158]= -834157373;
assign addr[18159]= -763158411;
assign addr[18160]= -691191324;
assign addr[18161]= -618347408;
assign addr[18162]= -544719071;
assign addr[18163]= -470399716;
assign addr[18164]= -395483624;
assign addr[18165]= -320065829;
assign addr[18166]= -244242007;
assign addr[18167]= -168108346;
assign addr[18168]= -91761426;
assign addr[18169]= -15298099;
assign addr[18170]= 61184634;
assign addr[18171]= 137589750;
assign addr[18172]= 213820322;
assign addr[18173]= 289779648;
assign addr[18174]= 365371365;
assign addr[18175]= 440499581;
assign addr[18176]= 515068990;
assign addr[18177]= 588984994;
assign addr[18178]= 662153826;
assign addr[18179]= 734482665;
assign addr[18180]= 805879757;
assign addr[18181]= 876254528;
assign addr[18182]= 945517704;
assign addr[18183]= 1013581418;
assign addr[18184]= 1080359326;
assign addr[18185]= 1145766716;
assign addr[18186]= 1209720613;
assign addr[18187]= 1272139887;
assign addr[18188]= 1332945355;
assign addr[18189]= 1392059879;
assign addr[18190]= 1449408469;
assign addr[18191]= 1504918373;
assign addr[18192]= 1558519173;
assign addr[18193]= 1610142873;
assign addr[18194]= 1659723983;
assign addr[18195]= 1707199606;
assign addr[18196]= 1752509516;
assign addr[18197]= 1795596234;
assign addr[18198]= 1836405100;
assign addr[18199]= 1874884346;
assign addr[18200]= 1910985158;
assign addr[18201]= 1944661739;
assign addr[18202]= 1975871368;
assign addr[18203]= 2004574453;
assign addr[18204]= 2030734582;
assign addr[18205]= 2054318569;
assign addr[18206]= 2075296495;
assign addr[18207]= 2093641749;
assign addr[18208]= 2109331059;
assign addr[18209]= 2122344521;
assign addr[18210]= 2132665626;
assign addr[18211]= 2140281282;
assign addr[18212]= 2145181827;
assign addr[18213]= 2147361045;
assign addr[18214]= 2146816171;
assign addr[18215]= 2143547897;
assign addr[18216]= 2137560369;
assign addr[18217]= 2128861181;
assign addr[18218]= 2117461370;
assign addr[18219]= 2103375398;
assign addr[18220]= 2086621133;
assign addr[18221]= 2067219829;
assign addr[18222]= 2045196100;
assign addr[18223]= 2020577882;
assign addr[18224]= 1993396407;
assign addr[18225]= 1963686155;
assign addr[18226]= 1931484818;
assign addr[18227]= 1896833245;
assign addr[18228]= 1859775393;
assign addr[18229]= 1820358275;
assign addr[18230]= 1778631892;
assign addr[18231]= 1734649179;
assign addr[18232]= 1688465931;
assign addr[18233]= 1640140734;
assign addr[18234]= 1589734894;
assign addr[18235]= 1537312353;
assign addr[18236]= 1482939614;
assign addr[18237]= 1426685652;
assign addr[18238]= 1368621831;
assign addr[18239]= 1308821808;
assign addr[18240]= 1247361445;
assign addr[18241]= 1184318708;
assign addr[18242]= 1119773573;
assign addr[18243]= 1053807919;
assign addr[18244]= 986505429;
assign addr[18245]= 917951481;
assign addr[18246]= 848233042;
assign addr[18247]= 777438554;
assign addr[18248]= 705657826;
assign addr[18249]= 632981917;
assign addr[18250]= 559503022;
assign addr[18251]= 485314355;
assign addr[18252]= 410510029;
assign addr[18253]= 335184940;
assign addr[18254]= 259434643;
assign addr[18255]= 183355234;
assign addr[18256]= 107043224;
assign addr[18257]= 30595422;
assign addr[18258]= -45891193;
assign addr[18259]= -122319591;
assign addr[18260]= -198592817;
assign addr[18261]= -274614114;
assign addr[18262]= -350287041;
assign addr[18263]= -425515602;
assign addr[18264]= -500204365;
assign addr[18265]= -574258580;
assign addr[18266]= -647584304;
assign addr[18267]= -720088517;
assign addr[18268]= -791679244;
assign addr[18269]= -862265664;
assign addr[18270]= -931758235;
assign addr[18271]= -1000068799;
assign addr[18272]= -1067110699;
assign addr[18273]= -1132798888;
assign addr[18274]= -1197050035;
assign addr[18275]= -1259782632;
assign addr[18276]= -1320917099;
assign addr[18277]= -1380375881;
assign addr[18278]= -1438083551;
assign addr[18279]= -1493966902;
assign addr[18280]= -1547955041;
assign addr[18281]= -1599979481;
assign addr[18282]= -1649974225;
assign addr[18283]= -1697875851;
assign addr[18284]= -1743623590;
assign addr[18285]= -1787159411;
assign addr[18286]= -1828428082;
assign addr[18287]= -1867377253;
assign addr[18288]= -1903957513;
assign addr[18289]= -1938122457;
assign addr[18290]= -1969828744;
assign addr[18291]= -1999036154;
assign addr[18292]= -2025707632;
assign addr[18293]= -2049809346;
assign addr[18294]= -2071310720;
assign addr[18295]= -2090184478;
assign addr[18296]= -2106406677;
assign addr[18297]= -2119956737;
assign addr[18298]= -2130817471;
assign addr[18299]= -2138975100;
assign addr[18300]= -2144419275;
assign addr[18301]= -2147143090;
assign addr[18302]= -2147143090;
assign addr[18303]= -2144419275;
assign addr[18304]= -2138975100;
assign addr[18305]= -2130817471;
assign addr[18306]= -2119956737;
assign addr[18307]= -2106406677;
assign addr[18308]= -2090184478;
assign addr[18309]= -2071310720;
assign addr[18310]= -2049809346;
assign addr[18311]= -2025707632;
assign addr[18312]= -1999036154;
assign addr[18313]= -1969828744;
assign addr[18314]= -1938122457;
assign addr[18315]= -1903957513;
assign addr[18316]= -1867377253;
assign addr[18317]= -1828428082;
assign addr[18318]= -1787159411;
assign addr[18319]= -1743623590;
assign addr[18320]= -1697875851;
assign addr[18321]= -1649974225;
assign addr[18322]= -1599979481;
assign addr[18323]= -1547955041;
assign addr[18324]= -1493966902;
assign addr[18325]= -1438083551;
assign addr[18326]= -1380375881;
assign addr[18327]= -1320917099;
assign addr[18328]= -1259782632;
assign addr[18329]= -1197050035;
assign addr[18330]= -1132798888;
assign addr[18331]= -1067110699;
assign addr[18332]= -1000068799;
assign addr[18333]= -931758235;
assign addr[18334]= -862265664;
assign addr[18335]= -791679244;
assign addr[18336]= -720088517;
assign addr[18337]= -647584304;
assign addr[18338]= -574258580;
assign addr[18339]= -500204365;
assign addr[18340]= -425515602;
assign addr[18341]= -350287041;
assign addr[18342]= -274614114;
assign addr[18343]= -198592817;
assign addr[18344]= -122319591;
assign addr[18345]= -45891193;
assign addr[18346]= 30595422;
assign addr[18347]= 107043224;
assign addr[18348]= 183355234;
assign addr[18349]= 259434643;
assign addr[18350]= 335184940;
assign addr[18351]= 410510029;
assign addr[18352]= 485314355;
assign addr[18353]= 559503022;
assign addr[18354]= 632981917;
assign addr[18355]= 705657826;
assign addr[18356]= 777438554;
assign addr[18357]= 848233042;
assign addr[18358]= 917951481;
assign addr[18359]= 986505429;
assign addr[18360]= 1053807919;
assign addr[18361]= 1119773573;
assign addr[18362]= 1184318708;
assign addr[18363]= 1247361445;
assign addr[18364]= 1308821808;
assign addr[18365]= 1368621831;
assign addr[18366]= 1426685652;
assign addr[18367]= 1482939614;
assign addr[18368]= 1537312353;
assign addr[18369]= 1589734894;
assign addr[18370]= 1640140734;
assign addr[18371]= 1688465931;
assign addr[18372]= 1734649179;
assign addr[18373]= 1778631892;
assign addr[18374]= 1820358275;
assign addr[18375]= 1859775393;
assign addr[18376]= 1896833245;
assign addr[18377]= 1931484818;
assign addr[18378]= 1963686155;
assign addr[18379]= 1993396407;
assign addr[18380]= 2020577882;
assign addr[18381]= 2045196100;
assign addr[18382]= 2067219829;
assign addr[18383]= 2086621133;
assign addr[18384]= 2103375398;
assign addr[18385]= 2117461370;
assign addr[18386]= 2128861181;
assign addr[18387]= 2137560369;
assign addr[18388]= 2143547897;
assign addr[18389]= 2146816171;
assign addr[18390]= 2147361045;
assign addr[18391]= 2145181827;
assign addr[18392]= 2140281282;
assign addr[18393]= 2132665626;
assign addr[18394]= 2122344521;
assign addr[18395]= 2109331059;
assign addr[18396]= 2093641749;
assign addr[18397]= 2075296495;
assign addr[18398]= 2054318569;
assign addr[18399]= 2030734582;
assign addr[18400]= 2004574453;
assign addr[18401]= 1975871368;
assign addr[18402]= 1944661739;
assign addr[18403]= 1910985158;
assign addr[18404]= 1874884346;
assign addr[18405]= 1836405100;
assign addr[18406]= 1795596234;
assign addr[18407]= 1752509516;
assign addr[18408]= 1707199606;
assign addr[18409]= 1659723983;
assign addr[18410]= 1610142873;
assign addr[18411]= 1558519173;
assign addr[18412]= 1504918373;
assign addr[18413]= 1449408469;
assign addr[18414]= 1392059879;
assign addr[18415]= 1332945355;
assign addr[18416]= 1272139887;
assign addr[18417]= 1209720613;
assign addr[18418]= 1145766716;
assign addr[18419]= 1080359326;
assign addr[18420]= 1013581418;
assign addr[18421]= 945517704;
assign addr[18422]= 876254528;
assign addr[18423]= 805879757;
assign addr[18424]= 734482665;
assign addr[18425]= 662153826;
assign addr[18426]= 588984994;
assign addr[18427]= 515068990;
assign addr[18428]= 440499581;
assign addr[18429]= 365371365;
assign addr[18430]= 289779648;
assign addr[18431]= 213820322;
assign addr[18432]= 137589750;
assign addr[18433]= 61184634;
assign addr[18434]= -15298099;
assign addr[18435]= -91761426;
assign addr[18436]= -168108346;
assign addr[18437]= -244242007;
assign addr[18438]= -320065829;
assign addr[18439]= -395483624;
assign addr[18440]= -470399716;
assign addr[18441]= -544719071;
assign addr[18442]= -618347408;
assign addr[18443]= -691191324;
assign addr[18444]= -763158411;
assign addr[18445]= -834157373;
assign addr[18446]= -904098143;
assign addr[18447]= -972891995;
assign addr[18448]= -1040451659;
assign addr[18449]= -1106691431;
assign addr[18450]= -1171527280;
assign addr[18451]= -1234876957;
assign addr[18452]= -1296660098;
assign addr[18453]= -1356798326;
assign addr[18454]= -1415215352;
assign addr[18455]= -1471837070;
assign addr[18456]= -1526591649;
assign addr[18457]= -1579409630;
assign addr[18458]= -1630224009;
assign addr[18459]= -1678970324;
assign addr[18460]= -1725586737;
assign addr[18461]= -1770014111;
assign addr[18462]= -1812196087;
assign addr[18463]= -1852079154;
assign addr[18464]= -1889612716;
assign addr[18465]= -1924749160;
assign addr[18466]= -1957443913;
assign addr[18467]= -1987655498;
assign addr[18468]= -2015345591;
assign addr[18469]= -2040479063;
assign addr[18470]= -2063024031;
assign addr[18471]= -2082951896;
assign addr[18472]= -2100237377;
assign addr[18473]= -2114858546;
assign addr[18474]= -2126796855;
assign addr[18475]= -2136037160;
assign addr[18476]= -2142567738;
assign addr[18477]= -2146380306;
assign addr[18478]= -2147470025;
assign addr[18479]= -2145835515;
assign addr[18480]= -2141478848;
assign addr[18481]= -2134405552;
assign addr[18482]= -2124624598;
assign addr[18483]= -2112148396;
assign addr[18484]= -2096992772;
assign addr[18485]= -2079176953;
assign addr[18486]= -2058723538;
assign addr[18487]= -2035658475;
assign addr[18488]= -2010011024;
assign addr[18489]= -1981813720;
assign addr[18490]= -1951102334;
assign addr[18491]= -1917915825;
assign addr[18492]= -1882296293;
assign addr[18493]= -1844288924;
assign addr[18494]= -1803941934;
assign addr[18495]= -1761306505;
assign addr[18496]= -1716436725;
assign addr[18497]= -1669389513;
assign addr[18498]= -1620224553;
assign addr[18499]= -1569004214;
assign addr[18500]= -1515793473;
assign addr[18501]= -1460659832;
assign addr[18502]= -1403673233;
assign addr[18503]= -1344905966;
assign addr[18504]= -1284432584;
assign addr[18505]= -1222329801;
assign addr[18506]= -1158676398;
assign addr[18507]= -1093553126;
assign addr[18508]= -1027042599;
assign addr[18509]= -959229189;
assign addr[18510]= -890198924;
assign addr[18511]= -820039373;
assign addr[18512]= -748839539;
assign addr[18513]= -676689746;
assign addr[18514]= -603681519;
assign addr[18515]= -529907477;
assign addr[18516]= -455461206;
assign addr[18517]= -380437148;
assign addr[18518]= -304930476;
assign addr[18519]= -229036977;
assign addr[18520]= -152852926;
assign addr[18521]= -76474970;
assign addr[18522]= 0;
assign addr[18523]= 76474970;
assign addr[18524]= 152852926;
assign addr[18525]= 229036977;
assign addr[18526]= 304930476;
assign addr[18527]= 380437148;
assign addr[18528]= 455461206;
assign addr[18529]= 529907477;
assign addr[18530]= 603681519;
assign addr[18531]= 676689746;
assign addr[18532]= 748839539;
assign addr[18533]= 820039373;
assign addr[18534]= 890198924;
assign addr[18535]= 959229189;
assign addr[18536]= 1027042599;
assign addr[18537]= 1093553126;
assign addr[18538]= 1158676398;
assign addr[18539]= 1222329801;
assign addr[18540]= 1284432584;
assign addr[18541]= 1344905966;
assign addr[18542]= 1403673233;
assign addr[18543]= 1460659832;
assign addr[18544]= 1515793473;
assign addr[18545]= 1569004214;
assign addr[18546]= 1620224553;
assign addr[18547]= 1669389513;
assign addr[18548]= 1716436725;
assign addr[18549]= 1761306505;
assign addr[18550]= 1803941934;
assign addr[18551]= 1844288924;
assign addr[18552]= 1882296293;
assign addr[18553]= 1917915825;
assign addr[18554]= 1951102334;
assign addr[18555]= 1981813720;
assign addr[18556]= 2010011024;
assign addr[18557]= 2035658475;
assign addr[18558]= 2058723538;
assign addr[18559]= 2079176953;
assign addr[18560]= 2096992772;
assign addr[18561]= 2112148396;
assign addr[18562]= 2124624598;
assign addr[18563]= 2134405552;
assign addr[18564]= 2141478848;
assign addr[18565]= 2145835515;
assign addr[18566]= 2147470025;
assign addr[18567]= 2146380306;
assign addr[18568]= 2142567738;
assign addr[18569]= 2136037160;
assign addr[18570]= 2126796855;
assign addr[18571]= 2114858546;
assign addr[18572]= 2100237377;
assign addr[18573]= 2082951896;
assign addr[18574]= 2063024031;
assign addr[18575]= 2040479063;
assign addr[18576]= 2015345591;
assign addr[18577]= 1987655498;
assign addr[18578]= 1957443913;
assign addr[18579]= 1924749160;
assign addr[18580]= 1889612716;
assign addr[18581]= 1852079154;
assign addr[18582]= 1812196087;
assign addr[18583]= 1770014111;
assign addr[18584]= 1725586737;
assign addr[18585]= 1678970324;
assign addr[18586]= 1630224009;
assign addr[18587]= 1579409630;
assign addr[18588]= 1526591649;
assign addr[18589]= 1471837070;
assign addr[18590]= 1415215352;
assign addr[18591]= 1356798326;
assign addr[18592]= 1296660098;
assign addr[18593]= 1234876957;
assign addr[18594]= 1171527280;
assign addr[18595]= 1106691431;
assign addr[18596]= 1040451659;
assign addr[18597]= 972891995;
assign addr[18598]= 904098143;
assign addr[18599]= 834157373;
assign addr[18600]= 763158411;
assign addr[18601]= 691191324;
assign addr[18602]= 618347408;
assign addr[18603]= 544719071;
assign addr[18604]= 470399716;
assign addr[18605]= 395483624;
assign addr[18606]= 320065829;
assign addr[18607]= 244242007;
assign addr[18608]= 168108346;
assign addr[18609]= 91761426;
assign addr[18610]= 15298099;
assign addr[18611]= -61184634;
assign addr[18612]= -137589750;
assign addr[18613]= -213820322;
assign addr[18614]= -289779648;
assign addr[18615]= -365371365;
assign addr[18616]= -440499581;
assign addr[18617]= -515068990;
assign addr[18618]= -588984994;
assign addr[18619]= -662153826;
assign addr[18620]= -734482665;
assign addr[18621]= -805879757;
assign addr[18622]= -876254528;
assign addr[18623]= -945517704;
assign addr[18624]= -1013581418;
assign addr[18625]= -1080359326;
assign addr[18626]= -1145766716;
assign addr[18627]= -1209720613;
assign addr[18628]= -1272139887;
assign addr[18629]= -1332945355;
assign addr[18630]= -1392059879;
assign addr[18631]= -1449408469;
assign addr[18632]= -1504918373;
assign addr[18633]= -1558519173;
assign addr[18634]= -1610142873;
assign addr[18635]= -1659723983;
assign addr[18636]= -1707199606;
assign addr[18637]= -1752509516;
assign addr[18638]= -1795596234;
assign addr[18639]= -1836405100;
assign addr[18640]= -1874884346;
assign addr[18641]= -1910985158;
assign addr[18642]= -1944661739;
assign addr[18643]= -1975871368;
assign addr[18644]= -2004574453;
assign addr[18645]= -2030734582;
assign addr[18646]= -2054318569;
assign addr[18647]= -2075296495;
assign addr[18648]= -2093641749;
assign addr[18649]= -2109331059;
assign addr[18650]= -2122344521;
assign addr[18651]= -2132665626;
assign addr[18652]= -2140281282;
assign addr[18653]= -2145181827;
assign addr[18654]= -2147361045;
assign addr[18655]= -2146816171;
assign addr[18656]= -2143547897;
assign addr[18657]= -2137560369;
assign addr[18658]= -2128861181;
assign addr[18659]= -2117461370;
assign addr[18660]= -2103375398;
assign addr[18661]= -2086621133;
assign addr[18662]= -2067219829;
assign addr[18663]= -2045196100;
assign addr[18664]= -2020577882;
assign addr[18665]= -1993396407;
assign addr[18666]= -1963686155;
assign addr[18667]= -1931484818;
assign addr[18668]= -1896833245;
assign addr[18669]= -1859775393;
assign addr[18670]= -1820358275;
assign addr[18671]= -1778631892;
assign addr[18672]= -1734649179;
assign addr[18673]= -1688465931;
assign addr[18674]= -1640140734;
assign addr[18675]= -1589734894;
assign addr[18676]= -1537312353;
assign addr[18677]= -1482939614;
assign addr[18678]= -1426685652;
assign addr[18679]= -1368621831;
assign addr[18680]= -1308821808;
assign addr[18681]= -1247361445;
assign addr[18682]= -1184318708;
assign addr[18683]= -1119773573;
assign addr[18684]= -1053807919;
assign addr[18685]= -986505429;
assign addr[18686]= -917951481;
assign addr[18687]= -848233042;
assign addr[18688]= -777438554;
assign addr[18689]= -705657826;
assign addr[18690]= -632981917;
assign addr[18691]= -559503022;
assign addr[18692]= -485314355;
assign addr[18693]= -410510029;
assign addr[18694]= -335184940;
assign addr[18695]= -259434643;
assign addr[18696]= -183355234;
assign addr[18697]= -107043224;
assign addr[18698]= -30595422;
assign addr[18699]= 45891193;
assign addr[18700]= 122319591;
assign addr[18701]= 198592817;
assign addr[18702]= 274614114;
assign addr[18703]= 350287041;
assign addr[18704]= 425515602;
assign addr[18705]= 500204365;
assign addr[18706]= 574258580;
assign addr[18707]= 647584304;
assign addr[18708]= 720088517;
assign addr[18709]= 791679244;
assign addr[18710]= 862265664;
assign addr[18711]= 931758235;
assign addr[18712]= 1000068799;
assign addr[18713]= 1067110699;
assign addr[18714]= 1132798888;
assign addr[18715]= 1197050035;
assign addr[18716]= 1259782632;
assign addr[18717]= 1320917099;
assign addr[18718]= 1380375881;
assign addr[18719]= 1438083551;
assign addr[18720]= 1493966902;
assign addr[18721]= 1547955041;
assign addr[18722]= 1599979481;
assign addr[18723]= 1649974225;
assign addr[18724]= 1697875851;
assign addr[18725]= 1743623590;
assign addr[18726]= 1787159411;
assign addr[18727]= 1828428082;
assign addr[18728]= 1867377253;
assign addr[18729]= 1903957513;
assign addr[18730]= 1938122457;
assign addr[18731]= 1969828744;
assign addr[18732]= 1999036154;
assign addr[18733]= 2025707632;
assign addr[18734]= 2049809346;
assign addr[18735]= 2071310720;
assign addr[18736]= 2090184478;
assign addr[18737]= 2106406677;
assign addr[18738]= 2119956737;
assign addr[18739]= 2130817471;
assign addr[18740]= 2138975100;
assign addr[18741]= 2144419275;
assign addr[18742]= 2147143090;
assign addr[18743]= 2147143090;
assign addr[18744]= 2144419275;
assign addr[18745]= 2138975100;
assign addr[18746]= 2130817471;
assign addr[18747]= 2119956737;
assign addr[18748]= 2106406677;
assign addr[18749]= 2090184478;
assign addr[18750]= 2071310720;
assign addr[18751]= 2049809346;
assign addr[18752]= 2025707632;
assign addr[18753]= 1999036154;
assign addr[18754]= 1969828744;
assign addr[18755]= 1938122457;
assign addr[18756]= 1903957513;
assign addr[18757]= 1867377253;
assign addr[18758]= 1828428082;
assign addr[18759]= 1787159411;
assign addr[18760]= 1743623590;
assign addr[18761]= 1697875851;
assign addr[18762]= 1649974225;
assign addr[18763]= 1599979481;
assign addr[18764]= 1547955041;
assign addr[18765]= 1493966902;
assign addr[18766]= 1438083551;
assign addr[18767]= 1380375881;
assign addr[18768]= 1320917099;
assign addr[18769]= 1259782632;
assign addr[18770]= 1197050035;
assign addr[18771]= 1132798888;
assign addr[18772]= 1067110699;
assign addr[18773]= 1000068799;
assign addr[18774]= 931758235;
assign addr[18775]= 862265664;
assign addr[18776]= 791679244;
assign addr[18777]= 720088517;
assign addr[18778]= 647584304;
assign addr[18779]= 574258580;
assign addr[18780]= 500204365;
assign addr[18781]= 425515602;
assign addr[18782]= 350287041;
assign addr[18783]= 274614114;
assign addr[18784]= 198592817;
assign addr[18785]= 122319591;
assign addr[18786]= 45891193;
assign addr[18787]= -30595422;
assign addr[18788]= -107043224;
assign addr[18789]= -183355234;
assign addr[18790]= -259434643;
assign addr[18791]= -335184940;
assign addr[18792]= -410510029;
assign addr[18793]= -485314355;
assign addr[18794]= -559503022;
assign addr[18795]= -632981917;
assign addr[18796]= -705657826;
assign addr[18797]= -777438554;
assign addr[18798]= -848233042;
assign addr[18799]= -917951481;
assign addr[18800]= -986505429;
assign addr[18801]= -1053807919;
assign addr[18802]= -1119773573;
assign addr[18803]= -1184318708;
assign addr[18804]= -1247361445;
assign addr[18805]= -1308821808;
assign addr[18806]= -1368621831;
assign addr[18807]= -1426685652;
assign addr[18808]= -1482939614;
assign addr[18809]= -1537312353;
assign addr[18810]= -1589734894;
assign addr[18811]= -1640140734;
assign addr[18812]= -1688465931;
assign addr[18813]= -1734649179;
assign addr[18814]= -1778631892;
assign addr[18815]= -1820358275;
assign addr[18816]= -1859775393;
assign addr[18817]= -1896833245;
assign addr[18818]= -1931484818;
assign addr[18819]= -1963686155;
assign addr[18820]= -1993396407;
assign addr[18821]= -2020577882;
assign addr[18822]= -2045196100;
assign addr[18823]= -2067219829;
assign addr[18824]= -2086621133;
assign addr[18825]= -2103375398;
assign addr[18826]= -2117461370;
assign addr[18827]= -2128861181;
assign addr[18828]= -2137560369;
assign addr[18829]= -2143547897;
assign addr[18830]= -2146816171;
assign addr[18831]= -2147361045;
assign addr[18832]= -2145181827;
assign addr[18833]= -2140281282;
assign addr[18834]= -2132665626;
assign addr[18835]= -2122344521;
assign addr[18836]= -2109331059;
assign addr[18837]= -2093641749;
assign addr[18838]= -2075296495;
assign addr[18839]= -2054318569;
assign addr[18840]= -2030734582;
assign addr[18841]= -2004574453;
assign addr[18842]= -1975871368;
assign addr[18843]= -1944661739;
assign addr[18844]= -1910985158;
assign addr[18845]= -1874884346;
assign addr[18846]= -1836405100;
assign addr[18847]= -1795596234;
assign addr[18848]= -1752509516;
assign addr[18849]= -1707199606;
assign addr[18850]= -1659723983;
assign addr[18851]= -1610142873;
assign addr[18852]= -1558519173;
assign addr[18853]= -1504918373;
assign addr[18854]= -1449408469;
assign addr[18855]= -1392059879;
assign addr[18856]= -1332945355;
assign addr[18857]= -1272139887;
assign addr[18858]= -1209720613;
assign addr[18859]= -1145766716;
assign addr[18860]= -1080359326;
assign addr[18861]= -1013581418;
assign addr[18862]= -945517704;
assign addr[18863]= -876254528;
assign addr[18864]= -805879757;
assign addr[18865]= -734482665;
assign addr[18866]= -662153826;
assign addr[18867]= -588984994;
assign addr[18868]= -515068990;
assign addr[18869]= -440499581;
assign addr[18870]= -365371365;
assign addr[18871]= -289779648;
assign addr[18872]= -213820322;
assign addr[18873]= -137589750;
assign addr[18874]= -61184634;
assign addr[18875]= 15298099;
assign addr[18876]= 91761426;
assign addr[18877]= 168108346;
assign addr[18878]= 244242007;
assign addr[18879]= 320065829;
assign addr[18880]= 395483624;
assign addr[18881]= 470399716;
assign addr[18882]= 544719071;
assign addr[18883]= 618347408;
assign addr[18884]= 691191324;
assign addr[18885]= 763158411;
assign addr[18886]= 834157373;
assign addr[18887]= 904098143;
assign addr[18888]= 972891995;
assign addr[18889]= 1040451659;
assign addr[18890]= 1106691431;
assign addr[18891]= 1171527280;
assign addr[18892]= 1234876957;
assign addr[18893]= 1296660098;
assign addr[18894]= 1356798326;
assign addr[18895]= 1415215352;
assign addr[18896]= 1471837070;
assign addr[18897]= 1526591649;
assign addr[18898]= 1579409630;
assign addr[18899]= 1630224009;
assign addr[18900]= 1678970324;
assign addr[18901]= 1725586737;
assign addr[18902]= 1770014111;
assign addr[18903]= 1812196087;
assign addr[18904]= 1852079154;
assign addr[18905]= 1889612716;
assign addr[18906]= 1924749160;
assign addr[18907]= 1957443913;
assign addr[18908]= 1987655498;
assign addr[18909]= 2015345591;
assign addr[18910]= 2040479063;
assign addr[18911]= 2063024031;
assign addr[18912]= 2082951896;
assign addr[18913]= 2100237377;
assign addr[18914]= 2114858546;
assign addr[18915]= 2126796855;
assign addr[18916]= 2136037160;
assign addr[18917]= 2142567738;
assign addr[18918]= 2146380306;
assign addr[18919]= 2147470025;
assign addr[18920]= 2145835515;
assign addr[18921]= 2141478848;
assign addr[18922]= 2134405552;
assign addr[18923]= 2124624598;
assign addr[18924]= 2112148396;
assign addr[18925]= 2096992772;
assign addr[18926]= 2079176953;
assign addr[18927]= 2058723538;
assign addr[18928]= 2035658475;
assign addr[18929]= 2010011024;
assign addr[18930]= 1981813720;
assign addr[18931]= 1951102334;
assign addr[18932]= 1917915825;
assign addr[18933]= 1882296293;
assign addr[18934]= 1844288924;
assign addr[18935]= 1803941934;
assign addr[18936]= 1761306505;
assign addr[18937]= 1716436725;
assign addr[18938]= 1669389513;
assign addr[18939]= 1620224553;
assign addr[18940]= 1569004214;
assign addr[18941]= 1515793473;
assign addr[18942]= 1460659832;
assign addr[18943]= 1403673233;
assign addr[18944]= 1344905966;
assign addr[18945]= 1284432584;
assign addr[18946]= 1222329801;
assign addr[18947]= 1158676398;
assign addr[18948]= 1093553126;
assign addr[18949]= 1027042599;
assign addr[18950]= 959229189;
assign addr[18951]= 890198924;
assign addr[18952]= 820039373;
assign addr[18953]= 748839539;
assign addr[18954]= 676689746;
assign addr[18955]= 603681519;
assign addr[18956]= 529907477;
assign addr[18957]= 455461206;
assign addr[18958]= 380437148;
assign addr[18959]= 304930476;
assign addr[18960]= 229036977;
assign addr[18961]= 152852926;
assign addr[18962]= 76474970;
assign addr[18963]= 0;
assign addr[18964]= -76474970;
assign addr[18965]= -152852926;
assign addr[18966]= -229036977;
assign addr[18967]= -304930476;
assign addr[18968]= -380437148;
assign addr[18969]= -455461206;
assign addr[18970]= -529907477;
assign addr[18971]= -603681519;
assign addr[18972]= -676689746;
assign addr[18973]= -748839539;
assign addr[18974]= -820039373;
assign addr[18975]= -890198924;
assign addr[18976]= -959229189;
assign addr[18977]= -1027042599;
assign addr[18978]= -1093553126;
assign addr[18979]= -1158676398;
assign addr[18980]= -1222329801;
assign addr[18981]= -1284432584;
assign addr[18982]= -1344905966;
assign addr[18983]= -1403673233;
assign addr[18984]= -1460659832;
assign addr[18985]= -1515793473;
assign addr[18986]= -1569004214;
assign addr[18987]= -1620224553;
assign addr[18988]= -1669389513;
assign addr[18989]= -1716436725;
assign addr[18990]= -1761306505;
assign addr[18991]= -1803941934;
assign addr[18992]= -1844288924;
assign addr[18993]= -1882296293;
assign addr[18994]= -1917915825;
assign addr[18995]= -1951102334;
assign addr[18996]= -1981813720;
assign addr[18997]= -2010011024;
assign addr[18998]= -2035658475;
assign addr[18999]= -2058723538;
assign addr[19000]= -2079176953;
assign addr[19001]= -2096992772;
assign addr[19002]= -2112148396;
assign addr[19003]= -2124624598;
assign addr[19004]= -2134405552;
assign addr[19005]= -2141478848;
assign addr[19006]= -2145835515;
assign addr[19007]= -2147470025;
assign addr[19008]= -2146380306;
assign addr[19009]= -2142567738;
assign addr[19010]= -2136037160;
assign addr[19011]= -2126796855;
assign addr[19012]= -2114858546;
assign addr[19013]= -2100237377;
assign addr[19014]= -2082951896;
assign addr[19015]= -2063024031;
assign addr[19016]= -2040479063;
assign addr[19017]= -2015345591;
assign addr[19018]= -1987655498;
assign addr[19019]= -1957443913;
assign addr[19020]= -1924749160;
assign addr[19021]= -1889612716;
assign addr[19022]= -1852079154;
assign addr[19023]= -1812196087;
assign addr[19024]= -1770014111;
assign addr[19025]= -1725586737;
assign addr[19026]= -1678970324;
assign addr[19027]= -1630224009;
assign addr[19028]= -1579409630;
assign addr[19029]= -1526591649;
assign addr[19030]= -1471837070;
assign addr[19031]= -1415215352;
assign addr[19032]= -1356798326;
assign addr[19033]= -1296660098;
assign addr[19034]= -1234876957;
assign addr[19035]= -1171527280;
assign addr[19036]= -1106691431;
assign addr[19037]= -1040451659;
assign addr[19038]= -972891995;
assign addr[19039]= -904098143;
assign addr[19040]= -834157373;
assign addr[19041]= -763158411;
assign addr[19042]= -691191324;
assign addr[19043]= -618347408;
assign addr[19044]= -544719071;
assign addr[19045]= -470399716;
assign addr[19046]= -395483624;
assign addr[19047]= -320065829;
assign addr[19048]= -244242007;
assign addr[19049]= -168108346;
assign addr[19050]= -91761426;
assign addr[19051]= -15298099;
assign addr[19052]= 61184634;
assign addr[19053]= 137589750;
assign addr[19054]= 213820322;
assign addr[19055]= 289779648;
assign addr[19056]= 365371365;
assign addr[19057]= 440499581;
assign addr[19058]= 515068990;
assign addr[19059]= 588984994;
assign addr[19060]= 662153826;
assign addr[19061]= 734482665;
assign addr[19062]= 805879757;
assign addr[19063]= 876254528;
assign addr[19064]= 945517704;
assign addr[19065]= 1013581418;
assign addr[19066]= 1080359326;
assign addr[19067]= 1145766716;
assign addr[19068]= 1209720613;
assign addr[19069]= 1272139887;
assign addr[19070]= 1332945355;
assign addr[19071]= 1392059879;
assign addr[19072]= 1449408469;
assign addr[19073]= 1504918373;
assign addr[19074]= 1558519173;
assign addr[19075]= 1610142873;
assign addr[19076]= 1659723983;
assign addr[19077]= 1707199606;
assign addr[19078]= 1752509516;
assign addr[19079]= 1795596234;
assign addr[19080]= 1836405100;
assign addr[19081]= 1874884346;
assign addr[19082]= 1910985158;
assign addr[19083]= 1944661739;
assign addr[19084]= 1975871368;
assign addr[19085]= 2004574453;
assign addr[19086]= 2030734582;
assign addr[19087]= 2054318569;
assign addr[19088]= 2075296495;
assign addr[19089]= 2093641749;
assign addr[19090]= 2109331059;
assign addr[19091]= 2122344521;
assign addr[19092]= 2132665626;
assign addr[19093]= 2140281282;
assign addr[19094]= 2145181827;
assign addr[19095]= 2147361045;
assign addr[19096]= 2146816171;
assign addr[19097]= 2143547897;
assign addr[19098]= 2137560369;
assign addr[19099]= 2128861181;
assign addr[19100]= 2117461370;
assign addr[19101]= 2103375398;
assign addr[19102]= 2086621133;
assign addr[19103]= 2067219829;
assign addr[19104]= 2045196100;
assign addr[19105]= 2020577882;
assign addr[19106]= 1993396407;
assign addr[19107]= 1963686155;
assign addr[19108]= 1931484818;
assign addr[19109]= 1896833245;
assign addr[19110]= 1859775393;
assign addr[19111]= 1820358275;
assign addr[19112]= 1778631892;
assign addr[19113]= 1734649179;
assign addr[19114]= 1688465931;
assign addr[19115]= 1640140734;
assign addr[19116]= 1589734894;
assign addr[19117]= 1537312353;
assign addr[19118]= 1482939614;
assign addr[19119]= 1426685652;
assign addr[19120]= 1368621831;
assign addr[19121]= 1308821808;
assign addr[19122]= 1247361445;
assign addr[19123]= 1184318708;
assign addr[19124]= 1119773573;
assign addr[19125]= 1053807919;
assign addr[19126]= 986505429;
assign addr[19127]= 917951481;
assign addr[19128]= 848233042;
assign addr[19129]= 777438554;
assign addr[19130]= 705657826;
assign addr[19131]= 632981917;
assign addr[19132]= 559503022;
assign addr[19133]= 485314355;
assign addr[19134]= 410510029;
assign addr[19135]= 335184940;
assign addr[19136]= 259434643;
assign addr[19137]= 183355234;
assign addr[19138]= 107043224;
assign addr[19139]= 30595422;
assign addr[19140]= -45891193;
assign addr[19141]= -122319591;
assign addr[19142]= -198592817;
assign addr[19143]= -274614114;
assign addr[19144]= -350287041;
assign addr[19145]= -425515602;
assign addr[19146]= -500204365;
assign addr[19147]= -574258580;
assign addr[19148]= -647584304;
assign addr[19149]= -720088517;
assign addr[19150]= -791679244;
assign addr[19151]= -862265664;
assign addr[19152]= -931758235;
assign addr[19153]= -1000068799;
assign addr[19154]= -1067110699;
assign addr[19155]= -1132798888;
assign addr[19156]= -1197050035;
assign addr[19157]= -1259782632;
assign addr[19158]= -1320917099;
assign addr[19159]= -1380375881;
assign addr[19160]= -1438083551;
assign addr[19161]= -1493966902;
assign addr[19162]= -1547955041;
assign addr[19163]= -1599979481;
assign addr[19164]= -1649974225;
assign addr[19165]= -1697875851;
assign addr[19166]= -1743623590;
assign addr[19167]= -1787159411;
assign addr[19168]= -1828428082;
assign addr[19169]= -1867377253;
assign addr[19170]= -1903957513;
assign addr[19171]= -1938122457;
assign addr[19172]= -1969828744;
assign addr[19173]= -1999036154;
assign addr[19174]= -2025707632;
assign addr[19175]= -2049809346;
assign addr[19176]= -2071310720;
assign addr[19177]= -2090184478;
assign addr[19178]= -2106406677;
assign addr[19179]= -2119956737;
assign addr[19180]= -2130817471;
assign addr[19181]= -2138975100;
assign addr[19182]= -2144419275;
assign addr[19183]= -2147143090;
assign addr[19184]= -2147143090;
assign addr[19185]= -2144419275;
assign addr[19186]= -2138975100;
assign addr[19187]= -2130817471;
assign addr[19188]= -2119956737;
assign addr[19189]= -2106406677;
assign addr[19190]= -2090184478;
assign addr[19191]= -2071310720;
assign addr[19192]= -2049809346;
assign addr[19193]= -2025707632;
assign addr[19194]= -1999036154;
assign addr[19195]= -1969828744;
assign addr[19196]= -1938122457;
assign addr[19197]= -1903957513;
assign addr[19198]= -1867377253;
assign addr[19199]= -1828428082;
assign addr[19200]= -1787159411;
assign addr[19201]= -1743623590;
assign addr[19202]= -1697875851;
assign addr[19203]= -1649974225;
assign addr[19204]= -1599979481;
assign addr[19205]= -1547955041;
assign addr[19206]= -1493966902;
assign addr[19207]= -1438083551;
assign addr[19208]= -1380375881;
assign addr[19209]= -1320917099;
assign addr[19210]= -1259782632;
assign addr[19211]= -1197050035;
assign addr[19212]= -1132798888;
assign addr[19213]= -1067110699;
assign addr[19214]= -1000068799;
assign addr[19215]= -931758235;
assign addr[19216]= -862265664;
assign addr[19217]= -791679244;
assign addr[19218]= -720088517;
assign addr[19219]= -647584304;
assign addr[19220]= -574258580;
assign addr[19221]= -500204365;
assign addr[19222]= -425515602;
assign addr[19223]= -350287041;
assign addr[19224]= -274614114;
assign addr[19225]= -198592817;
assign addr[19226]= -122319591;
assign addr[19227]= -45891193;
assign addr[19228]= 30595422;
assign addr[19229]= 107043224;
assign addr[19230]= 183355234;
assign addr[19231]= 259434643;
assign addr[19232]= 335184940;
assign addr[19233]= 410510029;
assign addr[19234]= 485314355;
assign addr[19235]= 559503022;
assign addr[19236]= 632981917;
assign addr[19237]= 705657826;
assign addr[19238]= 777438554;
assign addr[19239]= 848233042;
assign addr[19240]= 917951481;
assign addr[19241]= 986505429;
assign addr[19242]= 1053807919;
assign addr[19243]= 1119773573;
assign addr[19244]= 1184318708;
assign addr[19245]= 1247361445;
assign addr[19246]= 1308821808;
assign addr[19247]= 1368621831;
assign addr[19248]= 1426685652;
assign addr[19249]= 1482939614;
assign addr[19250]= 1537312353;
assign addr[19251]= 1589734894;
assign addr[19252]= 1640140734;
assign addr[19253]= 1688465931;
assign addr[19254]= 1734649179;
assign addr[19255]= 1778631892;
assign addr[19256]= 1820358275;
assign addr[19257]= 1859775393;
assign addr[19258]= 1896833245;
assign addr[19259]= 1931484818;
assign addr[19260]= 1963686155;
assign addr[19261]= 1993396407;
assign addr[19262]= 2020577882;
assign addr[19263]= 2045196100;
assign addr[19264]= 2067219829;
assign addr[19265]= 2086621133;
assign addr[19266]= 2103375398;
assign addr[19267]= 2117461370;
assign addr[19268]= 2128861181;
assign addr[19269]= 2137560369;
assign addr[19270]= 2143547897;
assign addr[19271]= 2146816171;
assign addr[19272]= 2147361045;
assign addr[19273]= 2145181827;
assign addr[19274]= 2140281282;
assign addr[19275]= 2132665626;
assign addr[19276]= 2122344521;
assign addr[19277]= 2109331059;
assign addr[19278]= 2093641749;
assign addr[19279]= 2075296495;
assign addr[19280]= 2054318569;
assign addr[19281]= 2030734582;
assign addr[19282]= 2004574453;
assign addr[19283]= 1975871368;
assign addr[19284]= 1944661739;
assign addr[19285]= 1910985158;
assign addr[19286]= 1874884346;
assign addr[19287]= 1836405100;
assign addr[19288]= 1795596234;
assign addr[19289]= 1752509516;
assign addr[19290]= 1707199606;
assign addr[19291]= 1659723983;
assign addr[19292]= 1610142873;
assign addr[19293]= 1558519173;
assign addr[19294]= 1504918373;
assign addr[19295]= 1449408469;
assign addr[19296]= 1392059879;
assign addr[19297]= 1332945355;
assign addr[19298]= 1272139887;
assign addr[19299]= 1209720613;
assign addr[19300]= 1145766716;
assign addr[19301]= 1080359326;
assign addr[19302]= 1013581418;
assign addr[19303]= 945517704;
assign addr[19304]= 876254528;
assign addr[19305]= 805879757;
assign addr[19306]= 734482665;
assign addr[19307]= 662153826;
assign addr[19308]= 588984994;
assign addr[19309]= 515068990;
assign addr[19310]= 440499581;
assign addr[19311]= 365371365;
assign addr[19312]= 289779648;
assign addr[19313]= 213820322;
assign addr[19314]= 137589750;
assign addr[19315]= 61184634;
assign addr[19316]= -15298099;
assign addr[19317]= -91761426;
assign addr[19318]= -168108346;
assign addr[19319]= -244242007;
assign addr[19320]= -320065829;
assign addr[19321]= -395483624;
assign addr[19322]= -470399716;
assign addr[19323]= -544719071;
assign addr[19324]= -618347408;
assign addr[19325]= -691191324;
assign addr[19326]= -763158411;
assign addr[19327]= -834157373;
assign addr[19328]= -904098143;
assign addr[19329]= -972891995;
assign addr[19330]= -1040451659;
assign addr[19331]= -1106691431;
assign addr[19332]= -1171527280;
assign addr[19333]= -1234876957;
assign addr[19334]= -1296660098;
assign addr[19335]= -1356798326;
assign addr[19336]= -1415215352;
assign addr[19337]= -1471837070;
assign addr[19338]= -1526591649;
assign addr[19339]= -1579409630;
assign addr[19340]= -1630224009;
assign addr[19341]= -1678970324;
assign addr[19342]= -1725586737;
assign addr[19343]= -1770014111;
assign addr[19344]= -1812196087;
assign addr[19345]= -1852079154;
assign addr[19346]= -1889612716;
assign addr[19347]= -1924749160;
assign addr[19348]= -1957443913;
assign addr[19349]= -1987655498;
assign addr[19350]= -2015345591;
assign addr[19351]= -2040479063;
assign addr[19352]= -2063024031;
assign addr[19353]= -2082951896;
assign addr[19354]= -2100237377;
assign addr[19355]= -2114858546;
assign addr[19356]= -2126796855;
assign addr[19357]= -2136037160;
assign addr[19358]= -2142567738;
assign addr[19359]= -2146380306;
assign addr[19360]= -2147470025;
assign addr[19361]= -2145835515;
assign addr[19362]= -2141478848;
assign addr[19363]= -2134405552;
assign addr[19364]= -2124624598;
assign addr[19365]= -2112148396;
assign addr[19366]= -2096992772;
assign addr[19367]= -2079176953;
assign addr[19368]= -2058723538;
assign addr[19369]= -2035658475;
assign addr[19370]= -2010011024;
assign addr[19371]= -1981813720;
assign addr[19372]= -1951102334;
assign addr[19373]= -1917915825;
assign addr[19374]= -1882296293;
assign addr[19375]= -1844288924;
assign addr[19376]= -1803941934;
assign addr[19377]= -1761306505;
assign addr[19378]= -1716436725;
assign addr[19379]= -1669389513;
assign addr[19380]= -1620224553;
assign addr[19381]= -1569004214;
assign addr[19382]= -1515793473;
assign addr[19383]= -1460659832;
assign addr[19384]= -1403673233;
assign addr[19385]= -1344905966;
assign addr[19386]= -1284432584;
assign addr[19387]= -1222329801;
assign addr[19388]= -1158676398;
assign addr[19389]= -1093553126;
assign addr[19390]= -1027042599;
assign addr[19391]= -959229189;
assign addr[19392]= -890198924;
assign addr[19393]= -820039373;
assign addr[19394]= -748839539;
assign addr[19395]= -676689746;
assign addr[19396]= -603681519;
assign addr[19397]= -529907477;
assign addr[19398]= -455461206;
assign addr[19399]= -380437148;
assign addr[19400]= -304930476;
assign addr[19401]= -229036977;
assign addr[19402]= -152852926;
assign addr[19403]= -76474970;
assign addr[19404]= 0;
assign addr[19405]= 76474970;
assign addr[19406]= 152852926;
assign addr[19407]= 229036977;
assign addr[19408]= 304930476;
assign addr[19409]= 380437148;
assign addr[19410]= 455461206;
assign addr[19411]= 529907477;
assign addr[19412]= 603681519;
assign addr[19413]= 676689746;
assign addr[19414]= 748839539;
assign addr[19415]= 820039373;
assign addr[19416]= 890198924;
assign addr[19417]= 959229189;
assign addr[19418]= 1027042599;
assign addr[19419]= 1093553126;
assign addr[19420]= 1158676398;
assign addr[19421]= 1222329801;
assign addr[19422]= 1284432584;
assign addr[19423]= 1344905966;
assign addr[19424]= 1403673233;
assign addr[19425]= 1460659832;
assign addr[19426]= 1515793473;
assign addr[19427]= 1569004214;
assign addr[19428]= 1620224553;
assign addr[19429]= 1669389513;
assign addr[19430]= 1716436725;
assign addr[19431]= 1761306505;
assign addr[19432]= 1803941934;
assign addr[19433]= 1844288924;
assign addr[19434]= 1882296293;
assign addr[19435]= 1917915825;
assign addr[19436]= 1951102334;
assign addr[19437]= 1981813720;
assign addr[19438]= 2010011024;
assign addr[19439]= 2035658475;
assign addr[19440]= 2058723538;
assign addr[19441]= 2079176953;
assign addr[19442]= 2096992772;
assign addr[19443]= 2112148396;
assign addr[19444]= 2124624598;
assign addr[19445]= 2134405552;
assign addr[19446]= 2141478848;
assign addr[19447]= 2145835515;
assign addr[19448]= 2147470025;
assign addr[19449]= 2146380306;
assign addr[19450]= 2142567738;
assign addr[19451]= 2136037160;
assign addr[19452]= 2126796855;
assign addr[19453]= 2114858546;
assign addr[19454]= 2100237377;
assign addr[19455]= 2082951896;
assign addr[19456]= 2063024031;
assign addr[19457]= 2040479063;
assign addr[19458]= 2015345591;
assign addr[19459]= 1987655498;
assign addr[19460]= 1957443913;
assign addr[19461]= 1924749160;
assign addr[19462]= 1889612716;
assign addr[19463]= 1852079154;
assign addr[19464]= 1812196087;
assign addr[19465]= 1770014111;
assign addr[19466]= 1725586737;
assign addr[19467]= 1678970324;
assign addr[19468]= 1630224009;
assign addr[19469]= 1579409630;
assign addr[19470]= 1526591649;
assign addr[19471]= 1471837070;
assign addr[19472]= 1415215352;
assign addr[19473]= 1356798326;
assign addr[19474]= 1296660098;
assign addr[19475]= 1234876957;
assign addr[19476]= 1171527280;
assign addr[19477]= 1106691431;
assign addr[19478]= 1040451659;
assign addr[19479]= 972891995;
assign addr[19480]= 904098143;
assign addr[19481]= 834157373;
assign addr[19482]= 763158411;
assign addr[19483]= 691191324;
assign addr[19484]= 618347408;
assign addr[19485]= 544719071;
assign addr[19486]= 470399716;
assign addr[19487]= 395483624;
assign addr[19488]= 320065829;
assign addr[19489]= 244242007;
assign addr[19490]= 168108346;
assign addr[19491]= 91761426;
assign addr[19492]= 15298099;
assign addr[19493]= -61184634;
assign addr[19494]= -137589750;
assign addr[19495]= -213820322;
assign addr[19496]= -289779648;
assign addr[19497]= -365371365;
assign addr[19498]= -440499581;
assign addr[19499]= -515068990;
assign addr[19500]= -588984994;
assign addr[19501]= -662153826;
assign addr[19502]= -734482665;
assign addr[19503]= -805879757;
assign addr[19504]= -876254528;
assign addr[19505]= -945517704;
assign addr[19506]= -1013581418;
assign addr[19507]= -1080359326;
assign addr[19508]= -1145766716;
assign addr[19509]= -1209720613;
assign addr[19510]= -1272139887;
assign addr[19511]= -1332945355;
assign addr[19512]= -1392059879;
assign addr[19513]= -1449408469;
assign addr[19514]= -1504918373;
assign addr[19515]= -1558519173;
assign addr[19516]= -1610142873;
assign addr[19517]= -1659723983;
assign addr[19518]= -1707199606;
assign addr[19519]= -1752509516;
assign addr[19520]= -1795596234;
assign addr[19521]= -1836405100;
assign addr[19522]= -1874884346;
assign addr[19523]= -1910985158;
assign addr[19524]= -1944661739;
assign addr[19525]= -1975871368;
assign addr[19526]= -2004574453;
assign addr[19527]= -2030734582;
assign addr[19528]= -2054318569;
assign addr[19529]= -2075296495;
assign addr[19530]= -2093641749;
assign addr[19531]= -2109331059;
assign addr[19532]= -2122344521;
assign addr[19533]= -2132665626;
assign addr[19534]= -2140281282;
assign addr[19535]= -2145181827;
assign addr[19536]= -2147361045;
assign addr[19537]= -2146816171;
assign addr[19538]= -2143547897;
assign addr[19539]= -2137560369;
assign addr[19540]= -2128861181;
assign addr[19541]= -2117461370;
assign addr[19542]= -2103375398;
assign addr[19543]= -2086621133;
assign addr[19544]= -2067219829;
assign addr[19545]= -2045196100;
assign addr[19546]= -2020577882;
assign addr[19547]= -1993396407;
assign addr[19548]= -1963686155;
assign addr[19549]= -1931484818;
assign addr[19550]= -1896833245;
assign addr[19551]= -1859775393;
assign addr[19552]= -1820358275;
assign addr[19553]= -1778631892;
assign addr[19554]= -1734649179;
assign addr[19555]= -1688465931;
assign addr[19556]= -1640140734;
assign addr[19557]= -1589734894;
assign addr[19558]= -1537312353;
assign addr[19559]= -1482939614;
assign addr[19560]= -1426685652;
assign addr[19561]= -1368621831;
assign addr[19562]= -1308821808;
assign addr[19563]= -1247361445;
assign addr[19564]= -1184318708;
assign addr[19565]= -1119773573;
assign addr[19566]= -1053807919;
assign addr[19567]= -986505429;
assign addr[19568]= -917951481;
assign addr[19569]= -848233042;
assign addr[19570]= -777438554;
assign addr[19571]= -705657826;
assign addr[19572]= -632981917;
assign addr[19573]= -559503022;
assign addr[19574]= -485314355;
assign addr[19575]= -410510029;
assign addr[19576]= -335184940;
assign addr[19577]= -259434643;
assign addr[19578]= -183355234;
assign addr[19579]= -107043224;
assign addr[19580]= -30595422;
assign addr[19581]= 45891193;
assign addr[19582]= 122319591;
assign addr[19583]= 198592817;
assign addr[19584]= 274614114;
assign addr[19585]= 350287041;
assign addr[19586]= 425515602;
assign addr[19587]= 500204365;
assign addr[19588]= 574258580;
assign addr[19589]= 647584304;
assign addr[19590]= 720088517;
assign addr[19591]= 791679244;
assign addr[19592]= 862265664;
assign addr[19593]= 931758235;
assign addr[19594]= 1000068799;
assign addr[19595]= 1067110699;
assign addr[19596]= 1132798888;
assign addr[19597]= 1197050035;
assign addr[19598]= 1259782632;
assign addr[19599]= 1320917099;
assign addr[19600]= 1380375881;
assign addr[19601]= 1438083551;
assign addr[19602]= 1493966902;
assign addr[19603]= 1547955041;
assign addr[19604]= 1599979481;
assign addr[19605]= 1649974225;
assign addr[19606]= 1697875851;
assign addr[19607]= 1743623590;
assign addr[19608]= 1787159411;
assign addr[19609]= 1828428082;
assign addr[19610]= 1867377253;
assign addr[19611]= 1903957513;
assign addr[19612]= 1938122457;
assign addr[19613]= 1969828744;
assign addr[19614]= 1999036154;
assign addr[19615]= 2025707632;
assign addr[19616]= 2049809346;
assign addr[19617]= 2071310720;
assign addr[19618]= 2090184478;
assign addr[19619]= 2106406677;
assign addr[19620]= 2119956737;
assign addr[19621]= 2130817471;
assign addr[19622]= 2138975100;
assign addr[19623]= 2144419275;
assign addr[19624]= 2147143090;
assign addr[19625]= 2147143090;
assign addr[19626]= 2144419275;
assign addr[19627]= 2138975100;
assign addr[19628]= 2130817471;
assign addr[19629]= 2119956737;
assign addr[19630]= 2106406677;
assign addr[19631]= 2090184478;
assign addr[19632]= 2071310720;
assign addr[19633]= 2049809346;
assign addr[19634]= 2025707632;
assign addr[19635]= 1999036154;
assign addr[19636]= 1969828744;
assign addr[19637]= 1938122457;
assign addr[19638]= 1903957513;
assign addr[19639]= 1867377253;
assign addr[19640]= 1828428082;
assign addr[19641]= 1787159411;
assign addr[19642]= 1743623590;
assign addr[19643]= 1697875851;
assign addr[19644]= 1649974225;
assign addr[19645]= 1599979481;
assign addr[19646]= 1547955041;
assign addr[19647]= 1493966902;
assign addr[19648]= 1438083551;
assign addr[19649]= 1380375881;
assign addr[19650]= 1320917099;
assign addr[19651]= 1259782632;
assign addr[19652]= 1197050035;
assign addr[19653]= 1132798888;
assign addr[19654]= 1067110699;
assign addr[19655]= 1000068799;
assign addr[19656]= 931758235;
assign addr[19657]= 862265664;
assign addr[19658]= 791679244;
assign addr[19659]= 720088517;
assign addr[19660]= 647584304;
assign addr[19661]= 574258580;
assign addr[19662]= 500204365;
assign addr[19663]= 425515602;
assign addr[19664]= 350287041;
assign addr[19665]= 274614114;
assign addr[19666]= 198592817;
assign addr[19667]= 122319591;
assign addr[19668]= 45891193;
assign addr[19669]= -30595422;
assign addr[19670]= -107043224;
assign addr[19671]= -183355234;
assign addr[19672]= -259434643;
assign addr[19673]= -335184940;
assign addr[19674]= -410510029;
assign addr[19675]= -485314355;
assign addr[19676]= -559503022;
assign addr[19677]= -632981917;
assign addr[19678]= -705657826;
assign addr[19679]= -777438554;
assign addr[19680]= -848233042;
assign addr[19681]= -917951481;
assign addr[19682]= -986505429;
assign addr[19683]= -1053807919;
assign addr[19684]= -1119773573;
assign addr[19685]= -1184318708;
assign addr[19686]= -1247361445;
assign addr[19687]= -1308821808;
assign addr[19688]= -1368621831;
assign addr[19689]= -1426685652;
assign addr[19690]= -1482939614;
assign addr[19691]= -1537312353;
assign addr[19692]= -1589734894;
assign addr[19693]= -1640140734;
assign addr[19694]= -1688465931;
assign addr[19695]= -1734649179;
assign addr[19696]= -1778631892;
assign addr[19697]= -1820358275;
assign addr[19698]= -1859775393;
assign addr[19699]= -1896833245;
assign addr[19700]= -1931484818;
assign addr[19701]= -1963686155;
assign addr[19702]= -1993396407;
assign addr[19703]= -2020577882;
assign addr[19704]= -2045196100;
assign addr[19705]= -2067219829;
assign addr[19706]= -2086621133;
assign addr[19707]= -2103375398;
assign addr[19708]= -2117461370;
assign addr[19709]= -2128861181;
assign addr[19710]= -2137560369;
assign addr[19711]= -2143547897;
assign addr[19712]= -2146816171;
assign addr[19713]= -2147361045;
assign addr[19714]= -2145181827;
assign addr[19715]= -2140281282;
assign addr[19716]= -2132665626;
assign addr[19717]= -2122344521;
assign addr[19718]= -2109331059;
assign addr[19719]= -2093641749;
assign addr[19720]= -2075296495;
assign addr[19721]= -2054318569;
assign addr[19722]= -2030734582;
assign addr[19723]= -2004574453;
assign addr[19724]= -1975871368;
assign addr[19725]= -1944661739;
assign addr[19726]= -1910985158;
assign addr[19727]= -1874884346;
assign addr[19728]= -1836405100;
assign addr[19729]= -1795596234;
assign addr[19730]= -1752509516;
assign addr[19731]= -1707199606;
assign addr[19732]= -1659723983;
assign addr[19733]= -1610142873;
assign addr[19734]= -1558519173;
assign addr[19735]= -1504918373;
assign addr[19736]= -1449408469;
assign addr[19737]= -1392059879;
assign addr[19738]= -1332945355;
assign addr[19739]= -1272139887;
assign addr[19740]= -1209720613;
assign addr[19741]= -1145766716;
assign addr[19742]= -1080359326;
assign addr[19743]= -1013581418;
assign addr[19744]= -945517704;
assign addr[19745]= -876254528;
assign addr[19746]= -805879757;
assign addr[19747]= -734482665;
assign addr[19748]= -662153826;
assign addr[19749]= -588984994;
assign addr[19750]= -515068990;
assign addr[19751]= -440499581;
assign addr[19752]= -365371365;
assign addr[19753]= -289779648;
assign addr[19754]= -213820322;
assign addr[19755]= -137589750;
assign addr[19756]= -61184634;
assign addr[19757]= 15298099;
assign addr[19758]= 91761426;
assign addr[19759]= 168108346;
assign addr[19760]= 244242007;
assign addr[19761]= 320065829;
assign addr[19762]= 395483624;
assign addr[19763]= 470399716;
assign addr[19764]= 544719071;
assign addr[19765]= 618347408;
assign addr[19766]= 691191324;
assign addr[19767]= 763158411;
assign addr[19768]= 834157373;
assign addr[19769]= 904098143;
assign addr[19770]= 972891995;
assign addr[19771]= 1040451659;
assign addr[19772]= 1106691431;
assign addr[19773]= 1171527280;
assign addr[19774]= 1234876957;
assign addr[19775]= 1296660098;
assign addr[19776]= 1356798326;
assign addr[19777]= 1415215352;
assign addr[19778]= 1471837070;
assign addr[19779]= 1526591649;
assign addr[19780]= 1579409630;
assign addr[19781]= 1630224009;
assign addr[19782]= 1678970324;
assign addr[19783]= 1725586737;
assign addr[19784]= 1770014111;
assign addr[19785]= 1812196087;
assign addr[19786]= 1852079154;
assign addr[19787]= 1889612716;
assign addr[19788]= 1924749160;
assign addr[19789]= 1957443913;
assign addr[19790]= 1987655498;
assign addr[19791]= 2015345591;
assign addr[19792]= 2040479063;
assign addr[19793]= 2063024031;
assign addr[19794]= 2082951896;
assign addr[19795]= 2100237377;
assign addr[19796]= 2114858546;
assign addr[19797]= 2126796855;
assign addr[19798]= 2136037160;
assign addr[19799]= 2142567738;
assign addr[19800]= 2146380306;
assign addr[19801]= 2147470025;
assign addr[19802]= 2145835515;
assign addr[19803]= 2141478848;
assign addr[19804]= 2134405552;
assign addr[19805]= 2124624598;
assign addr[19806]= 2112148396;
assign addr[19807]= 2096992772;
assign addr[19808]= 2079176953;
assign addr[19809]= 2058723538;
assign addr[19810]= 2035658475;
assign addr[19811]= 2010011024;
assign addr[19812]= 1981813720;
assign addr[19813]= 1951102334;
assign addr[19814]= 1917915825;
assign addr[19815]= 1882296293;
assign addr[19816]= 1844288924;
assign addr[19817]= 1803941934;
assign addr[19818]= 1761306505;
assign addr[19819]= 1716436725;
assign addr[19820]= 1669389513;
assign addr[19821]= 1620224553;
assign addr[19822]= 1569004214;
assign addr[19823]= 1515793473;
assign addr[19824]= 1460659832;
assign addr[19825]= 1403673233;
assign addr[19826]= 1344905966;
assign addr[19827]= 1284432584;
assign addr[19828]= 1222329801;
assign addr[19829]= 1158676398;
assign addr[19830]= 1093553126;
assign addr[19831]= 1027042599;
assign addr[19832]= 959229189;
assign addr[19833]= 890198924;
assign addr[19834]= 820039373;
assign addr[19835]= 748839539;
assign addr[19836]= 676689746;
assign addr[19837]= 603681519;
assign addr[19838]= 529907477;
assign addr[19839]= 455461206;
assign addr[19840]= 380437148;
assign addr[19841]= 304930476;
assign addr[19842]= 229036977;
assign addr[19843]= 152852926;
assign addr[19844]= 76474970;
assign addr[19845]= 0;
assign addr[19846]= -76474970;
assign addr[19847]= -152852926;
assign addr[19848]= -229036977;
assign addr[19849]= -304930476;
assign addr[19850]= -380437148;
assign addr[19851]= -455461206;
assign addr[19852]= -529907477;
assign addr[19853]= -603681519;
assign addr[19854]= -676689746;
assign addr[19855]= -748839539;
assign addr[19856]= -820039373;
assign addr[19857]= -890198924;
assign addr[19858]= -959229189;
assign addr[19859]= -1027042599;
assign addr[19860]= -1093553126;
assign addr[19861]= -1158676398;
assign addr[19862]= -1222329801;
assign addr[19863]= -1284432584;
assign addr[19864]= -1344905966;
assign addr[19865]= -1403673233;
assign addr[19866]= -1460659832;
assign addr[19867]= -1515793473;
assign addr[19868]= -1569004214;
assign addr[19869]= -1620224553;
assign addr[19870]= -1669389513;
assign addr[19871]= -1716436725;
assign addr[19872]= -1761306505;
assign addr[19873]= -1803941934;
assign addr[19874]= -1844288924;
assign addr[19875]= -1882296293;
assign addr[19876]= -1917915825;
assign addr[19877]= -1951102334;
assign addr[19878]= -1981813720;
assign addr[19879]= -2010011024;
assign addr[19880]= -2035658475;
assign addr[19881]= -2058723538;
assign addr[19882]= -2079176953;
assign addr[19883]= -2096992772;
assign addr[19884]= -2112148396;
assign addr[19885]= -2124624598;
assign addr[19886]= -2134405552;
assign addr[19887]= -2141478848;
assign addr[19888]= -2145835515;
assign addr[19889]= -2147470025;
assign addr[19890]= -2146380306;
assign addr[19891]= -2142567738;
assign addr[19892]= -2136037160;
assign addr[19893]= -2126796855;
assign addr[19894]= -2114858546;
assign addr[19895]= -2100237377;
assign addr[19896]= -2082951896;
assign addr[19897]= -2063024031;
assign addr[19898]= -2040479063;
assign addr[19899]= -2015345591;
assign addr[19900]= -1987655498;
assign addr[19901]= -1957443913;
assign addr[19902]= -1924749160;
assign addr[19903]= -1889612716;
assign addr[19904]= -1852079154;
assign addr[19905]= -1812196087;
assign addr[19906]= -1770014111;
assign addr[19907]= -1725586737;
assign addr[19908]= -1678970324;
assign addr[19909]= -1630224009;
assign addr[19910]= -1579409630;
assign addr[19911]= -1526591649;
assign addr[19912]= -1471837070;
assign addr[19913]= -1415215352;
assign addr[19914]= -1356798326;
assign addr[19915]= -1296660098;
assign addr[19916]= -1234876957;
assign addr[19917]= -1171527280;
assign addr[19918]= -1106691431;
assign addr[19919]= -1040451659;
assign addr[19920]= -972891995;
assign addr[19921]= -904098143;
assign addr[19922]= -834157373;
assign addr[19923]= -763158411;
assign addr[19924]= -691191324;
assign addr[19925]= -618347408;
assign addr[19926]= -544719071;
assign addr[19927]= -470399716;
assign addr[19928]= -395483624;
assign addr[19929]= -320065829;
assign addr[19930]= -244242007;
assign addr[19931]= -168108346;
assign addr[19932]= -91761426;
assign addr[19933]= -15298099;
assign addr[19934]= 61184634;
assign addr[19935]= 137589750;
assign addr[19936]= 213820322;
assign addr[19937]= 289779648;
assign addr[19938]= 365371365;
assign addr[19939]= 440499581;
assign addr[19940]= 515068990;
assign addr[19941]= 588984994;
assign addr[19942]= 662153826;
assign addr[19943]= 734482665;
assign addr[19944]= 805879757;
assign addr[19945]= 876254528;
assign addr[19946]= 945517704;
assign addr[19947]= 1013581418;
assign addr[19948]= 1080359326;
assign addr[19949]= 1145766716;
assign addr[19950]= 1209720613;
assign addr[19951]= 1272139887;
assign addr[19952]= 1332945355;
assign addr[19953]= 1392059879;
assign addr[19954]= 1449408469;
assign addr[19955]= 1504918373;
assign addr[19956]= 1558519173;
assign addr[19957]= 1610142873;
assign addr[19958]= 1659723983;
assign addr[19959]= 1707199606;
assign addr[19960]= 1752509516;
assign addr[19961]= 1795596234;
assign addr[19962]= 1836405100;
assign addr[19963]= 1874884346;
assign addr[19964]= 1910985158;
assign addr[19965]= 1944661739;
assign addr[19966]= 1975871368;
assign addr[19967]= 2004574453;
assign addr[19968]= 2030734582;
assign addr[19969]= 2054318569;
assign addr[19970]= 2075296495;
assign addr[19971]= 2093641749;
assign addr[19972]= 2109331059;
assign addr[19973]= 2122344521;
assign addr[19974]= 2132665626;
assign addr[19975]= 2140281282;
assign addr[19976]= 2145181827;
assign addr[19977]= 2147361045;
assign addr[19978]= 2146816171;
assign addr[19979]= 2143547897;
assign addr[19980]= 2137560369;
assign addr[19981]= 2128861181;
assign addr[19982]= 2117461370;
assign addr[19983]= 2103375398;
assign addr[19984]= 2086621133;
assign addr[19985]= 2067219829;
assign addr[19986]= 2045196100;
assign addr[19987]= 2020577882;
assign addr[19988]= 1993396407;
assign addr[19989]= 1963686155;
assign addr[19990]= 1931484818;
assign addr[19991]= 1896833245;
assign addr[19992]= 1859775393;
assign addr[19993]= 1820358275;
assign addr[19994]= 1778631892;
assign addr[19995]= 1734649179;
assign addr[19996]= 1688465931;
assign addr[19997]= 1640140734;
assign addr[19998]= 1589734894;
assign addr[19999]= 1537312353;
assign addr[20000]= 1482939614;
assign addr[20001]= 1426685652;
assign addr[20002]= 1368621831;
assign addr[20003]= 1308821808;
assign addr[20004]= 1247361445;
assign addr[20005]= 1184318708;
assign addr[20006]= 1119773573;
assign addr[20007]= 1053807919;
assign addr[20008]= 986505429;
assign addr[20009]= 917951481;
assign addr[20010]= 848233042;
assign addr[20011]= 777438554;
assign addr[20012]= 705657826;
assign addr[20013]= 632981917;
assign addr[20014]= 559503022;
assign addr[20015]= 485314355;
assign addr[20016]= 410510029;
assign addr[20017]= 335184940;
assign addr[20018]= 259434643;
assign addr[20019]= 183355234;
assign addr[20020]= 107043224;
assign addr[20021]= 30595422;
assign addr[20022]= -45891193;
assign addr[20023]= -122319591;
assign addr[20024]= -198592817;
assign addr[20025]= -274614114;
assign addr[20026]= -350287041;
assign addr[20027]= -425515602;
assign addr[20028]= -500204365;
assign addr[20029]= -574258580;
assign addr[20030]= -647584304;
assign addr[20031]= -720088517;
assign addr[20032]= -791679244;
assign addr[20033]= -862265664;
assign addr[20034]= -931758235;
assign addr[20035]= -1000068799;
assign addr[20036]= -1067110699;
assign addr[20037]= -1132798888;
assign addr[20038]= -1197050035;
assign addr[20039]= -1259782632;
assign addr[20040]= -1320917099;
assign addr[20041]= -1380375881;
assign addr[20042]= -1438083551;
assign addr[20043]= -1493966902;
assign addr[20044]= -1547955041;
assign addr[20045]= -1599979481;
assign addr[20046]= -1649974225;
assign addr[20047]= -1697875851;
assign addr[20048]= -1743623590;
assign addr[20049]= -1787159411;
assign addr[20050]= -1828428082;
assign addr[20051]= -1867377253;
assign addr[20052]= -1903957513;
assign addr[20053]= -1938122457;
assign addr[20054]= -1969828744;
assign addr[20055]= -1999036154;
assign addr[20056]= -2025707632;
assign addr[20057]= -2049809346;
assign addr[20058]= -2071310720;
assign addr[20059]= -2090184478;
assign addr[20060]= -2106406677;
assign addr[20061]= -2119956737;
assign addr[20062]= -2130817471;
assign addr[20063]= -2138975100;
assign addr[20064]= -2144419275;
assign addr[20065]= -2147143090;
assign addr[20066]= -2147143090;
assign addr[20067]= -2144419275;
assign addr[20068]= -2138975100;
assign addr[20069]= -2130817471;
assign addr[20070]= -2119956737;
assign addr[20071]= -2106406677;
assign addr[20072]= -2090184478;
assign addr[20073]= -2071310720;
assign addr[20074]= -2049809346;
assign addr[20075]= -2025707632;
assign addr[20076]= -1999036154;
assign addr[20077]= -1969828744;
assign addr[20078]= -1938122457;
assign addr[20079]= -1903957513;
assign addr[20080]= -1867377253;
assign addr[20081]= -1828428082;
assign addr[20082]= -1787159411;
assign addr[20083]= -1743623590;
assign addr[20084]= -1697875851;
assign addr[20085]= -1649974225;
assign addr[20086]= -1599979481;
assign addr[20087]= -1547955041;
assign addr[20088]= -1493966902;
assign addr[20089]= -1438083551;
assign addr[20090]= -1380375881;
assign addr[20091]= -1320917099;
assign addr[20092]= -1259782632;
assign addr[20093]= -1197050035;
assign addr[20094]= -1132798888;
assign addr[20095]= -1067110699;
assign addr[20096]= -1000068799;
assign addr[20097]= -931758235;
assign addr[20098]= -862265664;
assign addr[20099]= -791679244;
assign addr[20100]= -720088517;
assign addr[20101]= -647584304;
assign addr[20102]= -574258580;
assign addr[20103]= -500204365;
assign addr[20104]= -425515602;
assign addr[20105]= -350287041;
assign addr[20106]= -274614114;
assign addr[20107]= -198592817;
assign addr[20108]= -122319591;
assign addr[20109]= -45891193;
assign addr[20110]= 30595422;
assign addr[20111]= 107043224;
assign addr[20112]= 183355234;
assign addr[20113]= 259434643;
assign addr[20114]= 335184940;
assign addr[20115]= 410510029;
assign addr[20116]= 485314355;
assign addr[20117]= 559503022;
assign addr[20118]= 632981917;
assign addr[20119]= 705657826;
assign addr[20120]= 777438554;
assign addr[20121]= 848233042;
assign addr[20122]= 917951481;
assign addr[20123]= 986505429;
assign addr[20124]= 1053807919;
assign addr[20125]= 1119773573;
assign addr[20126]= 1184318708;
assign addr[20127]= 1247361445;
assign addr[20128]= 1308821808;
assign addr[20129]= 1368621831;
assign addr[20130]= 1426685652;
assign addr[20131]= 1482939614;
assign addr[20132]= 1537312353;
assign addr[20133]= 1589734894;
assign addr[20134]= 1640140734;
assign addr[20135]= 1688465931;
assign addr[20136]= 1734649179;
assign addr[20137]= 1778631892;
assign addr[20138]= 1820358275;
assign addr[20139]= 1859775393;
assign addr[20140]= 1896833245;
assign addr[20141]= 1931484818;
assign addr[20142]= 1963686155;
assign addr[20143]= 1993396407;
assign addr[20144]= 2020577882;
assign addr[20145]= 2045196100;
assign addr[20146]= 2067219829;
assign addr[20147]= 2086621133;
assign addr[20148]= 2103375398;
assign addr[20149]= 2117461370;
assign addr[20150]= 2128861181;
assign addr[20151]= 2137560369;
assign addr[20152]= 2143547897;
assign addr[20153]= 2146816171;
assign addr[20154]= 2147361045;
assign addr[20155]= 2145181827;
assign addr[20156]= 2140281282;
assign addr[20157]= 2132665626;
assign addr[20158]= 2122344521;
assign addr[20159]= 2109331059;
assign addr[20160]= 2093641749;
assign addr[20161]= 2075296495;
assign addr[20162]= 2054318569;
assign addr[20163]= 2030734582;
assign addr[20164]= 2004574453;
assign addr[20165]= 1975871368;
assign addr[20166]= 1944661739;
assign addr[20167]= 1910985158;
assign addr[20168]= 1874884346;
assign addr[20169]= 1836405100;
assign addr[20170]= 1795596234;
assign addr[20171]= 1752509516;
assign addr[20172]= 1707199606;
assign addr[20173]= 1659723983;
assign addr[20174]= 1610142873;
assign addr[20175]= 1558519173;
assign addr[20176]= 1504918373;
assign addr[20177]= 1449408469;
assign addr[20178]= 1392059879;
assign addr[20179]= 1332945355;
assign addr[20180]= 1272139887;
assign addr[20181]= 1209720613;
assign addr[20182]= 1145766716;
assign addr[20183]= 1080359326;
assign addr[20184]= 1013581418;
assign addr[20185]= 945517704;
assign addr[20186]= 876254528;
assign addr[20187]= 805879757;
assign addr[20188]= 734482665;
assign addr[20189]= 662153826;
assign addr[20190]= 588984994;
assign addr[20191]= 515068990;
assign addr[20192]= 440499581;
assign addr[20193]= 365371365;
assign addr[20194]= 289779648;
assign addr[20195]= 213820322;
assign addr[20196]= 137589750;
assign addr[20197]= 61184634;
assign addr[20198]= -15298099;
assign addr[20199]= -91761426;
assign addr[20200]= -168108346;
assign addr[20201]= -244242007;
assign addr[20202]= -320065829;
assign addr[20203]= -395483624;
assign addr[20204]= -470399716;
assign addr[20205]= -544719071;
assign addr[20206]= -618347408;
assign addr[20207]= -691191324;
assign addr[20208]= -763158411;
assign addr[20209]= -834157373;
assign addr[20210]= -904098143;
assign addr[20211]= -972891995;
assign addr[20212]= -1040451659;
assign addr[20213]= -1106691431;
assign addr[20214]= -1171527280;
assign addr[20215]= -1234876957;
assign addr[20216]= -1296660098;
assign addr[20217]= -1356798326;
assign addr[20218]= -1415215352;
assign addr[20219]= -1471837070;
assign addr[20220]= -1526591649;
assign addr[20221]= -1579409630;
assign addr[20222]= -1630224009;
assign addr[20223]= -1678970324;
assign addr[20224]= -1725586737;
assign addr[20225]= -1770014111;
assign addr[20226]= -1812196087;
assign addr[20227]= -1852079154;
assign addr[20228]= -1889612716;
assign addr[20229]= -1924749160;
assign addr[20230]= -1957443913;
assign addr[20231]= -1987655498;
assign addr[20232]= -2015345591;
assign addr[20233]= -2040479063;
assign addr[20234]= -2063024031;
assign addr[20235]= -2082951896;
assign addr[20236]= -2100237377;
assign addr[20237]= -2114858546;
assign addr[20238]= -2126796855;
assign addr[20239]= -2136037160;
assign addr[20240]= -2142567738;
assign addr[20241]= -2146380306;
assign addr[20242]= -2147470025;
assign addr[20243]= -2145835515;
assign addr[20244]= -2141478848;
assign addr[20245]= -2134405552;
assign addr[20246]= -2124624598;
assign addr[20247]= -2112148396;
assign addr[20248]= -2096992772;
assign addr[20249]= -2079176953;
assign addr[20250]= -2058723538;
assign addr[20251]= -2035658475;
assign addr[20252]= -2010011024;
assign addr[20253]= -1981813720;
assign addr[20254]= -1951102334;
assign addr[20255]= -1917915825;
assign addr[20256]= -1882296293;
assign addr[20257]= -1844288924;
assign addr[20258]= -1803941934;
assign addr[20259]= -1761306505;
assign addr[20260]= -1716436725;
assign addr[20261]= -1669389513;
assign addr[20262]= -1620224553;
assign addr[20263]= -1569004214;
assign addr[20264]= -1515793473;
assign addr[20265]= -1460659832;
assign addr[20266]= -1403673233;
assign addr[20267]= -1344905966;
assign addr[20268]= -1284432584;
assign addr[20269]= -1222329801;
assign addr[20270]= -1158676398;
assign addr[20271]= -1093553126;
assign addr[20272]= -1027042599;
assign addr[20273]= -959229189;
assign addr[20274]= -890198924;
assign addr[20275]= -820039373;
assign addr[20276]= -748839539;
assign addr[20277]= -676689746;
assign addr[20278]= -603681519;
assign addr[20279]= -529907477;
assign addr[20280]= -455461206;
assign addr[20281]= -380437148;
assign addr[20282]= -304930476;
assign addr[20283]= -229036977;
assign addr[20284]= -152852926;
assign addr[20285]= -76474970;
assign addr[20286]= 0;
assign addr[20287]= 76474970;
assign addr[20288]= 152852926;
assign addr[20289]= 229036977;
assign addr[20290]= 304930476;
assign addr[20291]= 380437148;
assign addr[20292]= 455461206;
assign addr[20293]= 529907477;
assign addr[20294]= 603681519;
assign addr[20295]= 676689746;
assign addr[20296]= 748839539;
assign addr[20297]= 820039373;
assign addr[20298]= 890198924;
assign addr[20299]= 959229189;
assign addr[20300]= 1027042599;
assign addr[20301]= 1093553126;
assign addr[20302]= 1158676398;
assign addr[20303]= 1222329801;
assign addr[20304]= 1284432584;
assign addr[20305]= 1344905966;
assign addr[20306]= 1403673233;
assign addr[20307]= 1460659832;
assign addr[20308]= 1515793473;
assign addr[20309]= 1569004214;
assign addr[20310]= 1620224553;
assign addr[20311]= 1669389513;
assign addr[20312]= 1716436725;
assign addr[20313]= 1761306505;
assign addr[20314]= 1803941934;
assign addr[20315]= 1844288924;
assign addr[20316]= 1882296293;
assign addr[20317]= 1917915825;
assign addr[20318]= 1951102334;
assign addr[20319]= 1981813720;
assign addr[20320]= 2010011024;
assign addr[20321]= 2035658475;
assign addr[20322]= 2058723538;
assign addr[20323]= 2079176953;
assign addr[20324]= 2096992772;
assign addr[20325]= 2112148396;
assign addr[20326]= 2124624598;
assign addr[20327]= 2134405552;
assign addr[20328]= 2141478848;
assign addr[20329]= 2145835515;
assign addr[20330]= 2147470025;
assign addr[20331]= 2146380306;
assign addr[20332]= 2142567738;
assign addr[20333]= 2136037160;
assign addr[20334]= 2126796855;
assign addr[20335]= 2114858546;
assign addr[20336]= 2100237377;
assign addr[20337]= 2082951896;
assign addr[20338]= 2063024031;
assign addr[20339]= 2040479063;
assign addr[20340]= 2015345591;
assign addr[20341]= 1987655498;
assign addr[20342]= 1957443913;
assign addr[20343]= 1924749160;
assign addr[20344]= 1889612716;
assign addr[20345]= 1852079154;
assign addr[20346]= 1812196087;
assign addr[20347]= 1770014111;
assign addr[20348]= 1725586737;
assign addr[20349]= 1678970324;
assign addr[20350]= 1630224009;
assign addr[20351]= 1579409630;
assign addr[20352]= 1526591649;
assign addr[20353]= 1471837070;
assign addr[20354]= 1415215352;
assign addr[20355]= 1356798326;
assign addr[20356]= 1296660098;
assign addr[20357]= 1234876957;
assign addr[20358]= 1171527280;
assign addr[20359]= 1106691431;
assign addr[20360]= 1040451659;
assign addr[20361]= 972891995;
assign addr[20362]= 904098143;
assign addr[20363]= 834157373;
assign addr[20364]= 763158411;
assign addr[20365]= 691191324;
assign addr[20366]= 618347408;
assign addr[20367]= 544719071;
assign addr[20368]= 470399716;
assign addr[20369]= 395483624;
assign addr[20370]= 320065829;
assign addr[20371]= 244242007;
assign addr[20372]= 168108346;
assign addr[20373]= 91761426;
assign addr[20374]= 15298099;
assign addr[20375]= -61184634;
assign addr[20376]= -137589750;
assign addr[20377]= -213820322;
assign addr[20378]= -289779648;
assign addr[20379]= -365371365;
assign addr[20380]= -440499581;
assign addr[20381]= -515068990;
assign addr[20382]= -588984994;
assign addr[20383]= -662153826;
assign addr[20384]= -734482665;
assign addr[20385]= -805879757;
assign addr[20386]= -876254528;
assign addr[20387]= -945517704;
assign addr[20388]= -1013581418;
assign addr[20389]= -1080359326;
assign addr[20390]= -1145766716;
assign addr[20391]= -1209720613;
assign addr[20392]= -1272139887;
assign addr[20393]= -1332945355;
assign addr[20394]= -1392059879;
assign addr[20395]= -1449408469;
assign addr[20396]= -1504918373;
assign addr[20397]= -1558519173;
assign addr[20398]= -1610142873;
assign addr[20399]= -1659723983;
assign addr[20400]= -1707199606;
assign addr[20401]= -1752509516;
assign addr[20402]= -1795596234;
assign addr[20403]= -1836405100;
assign addr[20404]= -1874884346;
assign addr[20405]= -1910985158;
assign addr[20406]= -1944661739;
assign addr[20407]= -1975871368;
assign addr[20408]= -2004574453;
assign addr[20409]= -2030734582;
assign addr[20410]= -2054318569;
assign addr[20411]= -2075296495;
assign addr[20412]= -2093641749;
assign addr[20413]= -2109331059;
assign addr[20414]= -2122344521;
assign addr[20415]= -2132665626;
assign addr[20416]= -2140281282;
assign addr[20417]= -2145181827;
assign addr[20418]= -2147361045;
assign addr[20419]= -2146816171;
assign addr[20420]= -2143547897;
assign addr[20421]= -2137560369;
assign addr[20422]= -2128861181;
assign addr[20423]= -2117461370;
assign addr[20424]= -2103375398;
assign addr[20425]= -2086621133;
assign addr[20426]= -2067219829;
assign addr[20427]= -2045196100;
assign addr[20428]= -2020577882;
assign addr[20429]= -1993396407;
assign addr[20430]= -1963686155;
assign addr[20431]= -1931484818;
assign addr[20432]= -1896833245;
assign addr[20433]= -1859775393;
assign addr[20434]= -1820358275;
assign addr[20435]= -1778631892;
assign addr[20436]= -1734649179;
assign addr[20437]= -1688465931;
assign addr[20438]= -1640140734;
assign addr[20439]= -1589734894;
assign addr[20440]= -1537312353;
assign addr[20441]= -1482939614;
assign addr[20442]= -1426685652;
assign addr[20443]= -1368621831;
assign addr[20444]= -1308821808;
assign addr[20445]= -1247361445;
assign addr[20446]= -1184318708;
assign addr[20447]= -1119773573;
assign addr[20448]= -1053807919;
assign addr[20449]= -986505429;
assign addr[20450]= -917951481;
assign addr[20451]= -848233042;
assign addr[20452]= -777438554;
assign addr[20453]= -705657826;
assign addr[20454]= -632981917;
assign addr[20455]= -559503022;
assign addr[20456]= -485314355;
assign addr[20457]= -410510029;
assign addr[20458]= -335184940;
assign addr[20459]= -259434643;
assign addr[20460]= -183355234;
assign addr[20461]= -107043224;
assign addr[20462]= -30595422;
assign addr[20463]= 45891193;
assign addr[20464]= 122319591;
assign addr[20465]= 198592817;
assign addr[20466]= 274614114;
assign addr[20467]= 350287041;
assign addr[20468]= 425515602;
assign addr[20469]= 500204365;
assign addr[20470]= 574258580;
assign addr[20471]= 647584304;
assign addr[20472]= 720088517;
assign addr[20473]= 791679244;
assign addr[20474]= 862265664;
assign addr[20475]= 931758235;
assign addr[20476]= 1000068799;
assign addr[20477]= 1067110699;
assign addr[20478]= 1132798888;
assign addr[20479]= 1197050035;
assign addr[20480]= 1259782632;
assign addr[20481]= 1320917099;
assign addr[20482]= 1380375881;
assign addr[20483]= 1438083551;
assign addr[20484]= 1493966902;
assign addr[20485]= 1547955041;
assign addr[20486]= 1599979481;
assign addr[20487]= 1649974225;
assign addr[20488]= 1697875851;
assign addr[20489]= 1743623590;
assign addr[20490]= 1787159411;
assign addr[20491]= 1828428082;
assign addr[20492]= 1867377253;
assign addr[20493]= 1903957513;
assign addr[20494]= 1938122457;
assign addr[20495]= 1969828744;
assign addr[20496]= 1999036154;
assign addr[20497]= 2025707632;
assign addr[20498]= 2049809346;
assign addr[20499]= 2071310720;
assign addr[20500]= 2090184478;
assign addr[20501]= 2106406677;
assign addr[20502]= 2119956737;
assign addr[20503]= 2130817471;
assign addr[20504]= 2138975100;
assign addr[20505]= 2144419275;
assign addr[20506]= 2147143090;
assign addr[20507]= 2147143090;
assign addr[20508]= 2144419275;
assign addr[20509]= 2138975100;
assign addr[20510]= 2130817471;
assign addr[20511]= 2119956737;
assign addr[20512]= 2106406677;
assign addr[20513]= 2090184478;
assign addr[20514]= 2071310720;
assign addr[20515]= 2049809346;
assign addr[20516]= 2025707632;
assign addr[20517]= 1999036154;
assign addr[20518]= 1969828744;
assign addr[20519]= 1938122457;
assign addr[20520]= 1903957513;
assign addr[20521]= 1867377253;
assign addr[20522]= 1828428082;
assign addr[20523]= 1787159411;
assign addr[20524]= 1743623590;
assign addr[20525]= 1697875851;
assign addr[20526]= 1649974225;
assign addr[20527]= 1599979481;
assign addr[20528]= 1547955041;
assign addr[20529]= 1493966902;
assign addr[20530]= 1438083551;
assign addr[20531]= 1380375881;
assign addr[20532]= 1320917099;
assign addr[20533]= 1259782632;
assign addr[20534]= 1197050035;
assign addr[20535]= 1132798888;
assign addr[20536]= 1067110699;
assign addr[20537]= 1000068799;
assign addr[20538]= 931758235;
assign addr[20539]= 862265664;
assign addr[20540]= 791679244;
assign addr[20541]= 720088517;
assign addr[20542]= 647584304;
assign addr[20543]= 574258580;
assign addr[20544]= 500204365;
assign addr[20545]= 425515602;
assign addr[20546]= 350287041;
assign addr[20547]= 274614114;
assign addr[20548]= 198592817;
assign addr[20549]= 122319591;
assign addr[20550]= 45891193;
assign addr[20551]= -30595422;
assign addr[20552]= -107043224;
assign addr[20553]= -183355234;
assign addr[20554]= -259434643;
assign addr[20555]= -335184940;
assign addr[20556]= -410510029;
assign addr[20557]= -485314355;
assign addr[20558]= -559503022;
assign addr[20559]= -632981917;
assign addr[20560]= -705657826;
assign addr[20561]= -777438554;
assign addr[20562]= -848233042;
assign addr[20563]= -917951481;
assign addr[20564]= -986505429;
assign addr[20565]= -1053807919;
assign addr[20566]= -1119773573;
assign addr[20567]= -1184318708;
assign addr[20568]= -1247361445;
assign addr[20569]= -1308821808;
assign addr[20570]= -1368621831;
assign addr[20571]= -1426685652;
assign addr[20572]= -1482939614;
assign addr[20573]= -1537312353;
assign addr[20574]= -1589734894;
assign addr[20575]= -1640140734;
assign addr[20576]= -1688465931;
assign addr[20577]= -1734649179;
assign addr[20578]= -1778631892;
assign addr[20579]= -1820358275;
assign addr[20580]= -1859775393;
assign addr[20581]= -1896833245;
assign addr[20582]= -1931484818;
assign addr[20583]= -1963686155;
assign addr[20584]= -1993396407;
assign addr[20585]= -2020577882;
assign addr[20586]= -2045196100;
assign addr[20587]= -2067219829;
assign addr[20588]= -2086621133;
assign addr[20589]= -2103375398;
assign addr[20590]= -2117461370;
assign addr[20591]= -2128861181;
assign addr[20592]= -2137560369;
assign addr[20593]= -2143547897;
assign addr[20594]= -2146816171;
assign addr[20595]= -2147361045;
assign addr[20596]= -2145181827;
assign addr[20597]= -2140281282;
assign addr[20598]= -2132665626;
assign addr[20599]= -2122344521;
assign addr[20600]= -2109331059;
assign addr[20601]= -2093641749;
assign addr[20602]= -2075296495;
assign addr[20603]= -2054318569;
assign addr[20604]= -2030734582;
assign addr[20605]= -2004574453;
assign addr[20606]= -1975871368;
assign addr[20607]= -1944661739;
assign addr[20608]= -1910985158;
assign addr[20609]= -1874884346;
assign addr[20610]= -1836405100;
assign addr[20611]= -1795596234;
assign addr[20612]= -1752509516;
assign addr[20613]= -1707199606;
assign addr[20614]= -1659723983;
assign addr[20615]= -1610142873;
assign addr[20616]= -1558519173;
assign addr[20617]= -1504918373;
assign addr[20618]= -1449408469;
assign addr[20619]= -1392059879;
assign addr[20620]= -1332945355;
assign addr[20621]= -1272139887;
assign addr[20622]= -1209720613;
assign addr[20623]= -1145766716;
assign addr[20624]= -1080359326;
assign addr[20625]= -1013581418;
assign addr[20626]= -945517704;
assign addr[20627]= -876254528;
assign addr[20628]= -805879757;
assign addr[20629]= -734482665;
assign addr[20630]= -662153826;
assign addr[20631]= -588984994;
assign addr[20632]= -515068990;
assign addr[20633]= -440499581;
assign addr[20634]= -365371365;
assign addr[20635]= -289779648;
assign addr[20636]= -213820322;
assign addr[20637]= -137589750;
assign addr[20638]= -61184634;
assign addr[20639]= 15298099;
assign addr[20640]= 91761426;
assign addr[20641]= 168108346;
assign addr[20642]= 244242007;
assign addr[20643]= 320065829;
assign addr[20644]= 395483624;
assign addr[20645]= 470399716;
assign addr[20646]= 544719071;
assign addr[20647]= 618347408;
assign addr[20648]= 691191324;
assign addr[20649]= 763158411;
assign addr[20650]= 834157373;
assign addr[20651]= 904098143;
assign addr[20652]= 972891995;
assign addr[20653]= 1040451659;
assign addr[20654]= 1106691431;
assign addr[20655]= 1171527280;
assign addr[20656]= 1234876957;
assign addr[20657]= 1296660098;
assign addr[20658]= 1356798326;
assign addr[20659]= 1415215352;
assign addr[20660]= 1471837070;
assign addr[20661]= 1526591649;
assign addr[20662]= 1579409630;
assign addr[20663]= 1630224009;
assign addr[20664]= 1678970324;
assign addr[20665]= 1725586737;
assign addr[20666]= 1770014111;
assign addr[20667]= 1812196087;
assign addr[20668]= 1852079154;
assign addr[20669]= 1889612716;
assign addr[20670]= 1924749160;
assign addr[20671]= 1957443913;
assign addr[20672]= 1987655498;
assign addr[20673]= 2015345591;
assign addr[20674]= 2040479063;
assign addr[20675]= 2063024031;
assign addr[20676]= 2082951896;
assign addr[20677]= 2100237377;
assign addr[20678]= 2114858546;
assign addr[20679]= 2126796855;
assign addr[20680]= 2136037160;
assign addr[20681]= 2142567738;
assign addr[20682]= 2146380306;
assign addr[20683]= 2147470025;
assign addr[20684]= 2145835515;
assign addr[20685]= 2141478848;
assign addr[20686]= 2134405552;
assign addr[20687]= 2124624598;
assign addr[20688]= 2112148396;
assign addr[20689]= 2096992772;
assign addr[20690]= 2079176953;
assign addr[20691]= 2058723538;
assign addr[20692]= 2035658475;
assign addr[20693]= 2010011024;
assign addr[20694]= 1981813720;
assign addr[20695]= 1951102334;
assign addr[20696]= 1917915825;
assign addr[20697]= 1882296293;
assign addr[20698]= 1844288924;
assign addr[20699]= 1803941934;
assign addr[20700]= 1761306505;
assign addr[20701]= 1716436725;
assign addr[20702]= 1669389513;
assign addr[20703]= 1620224553;
assign addr[20704]= 1569004214;
assign addr[20705]= 1515793473;
assign addr[20706]= 1460659832;
assign addr[20707]= 1403673233;
assign addr[20708]= 1344905966;
assign addr[20709]= 1284432584;
assign addr[20710]= 1222329801;
assign addr[20711]= 1158676398;
assign addr[20712]= 1093553126;
assign addr[20713]= 1027042599;
assign addr[20714]= 959229189;
assign addr[20715]= 890198924;
assign addr[20716]= 820039373;
assign addr[20717]= 748839539;
assign addr[20718]= 676689746;
assign addr[20719]= 603681519;
assign addr[20720]= 529907477;
assign addr[20721]= 455461206;
assign addr[20722]= 380437148;
assign addr[20723]= 304930476;
assign addr[20724]= 229036977;
assign addr[20725]= 152852926;
assign addr[20726]= 76474970;
assign addr[20727]= 0;
assign addr[20728]= -76474970;
assign addr[20729]= -152852926;
assign addr[20730]= -229036977;
assign addr[20731]= -304930476;
assign addr[20732]= -380437148;
assign addr[20733]= -455461206;
assign addr[20734]= -529907477;
assign addr[20735]= -603681519;
assign addr[20736]= -676689746;
assign addr[20737]= -748839539;
assign addr[20738]= -820039373;
assign addr[20739]= -890198924;
assign addr[20740]= -959229189;
assign addr[20741]= -1027042599;
assign addr[20742]= -1093553126;
assign addr[20743]= -1158676398;
assign addr[20744]= -1222329801;
assign addr[20745]= -1284432584;
assign addr[20746]= -1344905966;
assign addr[20747]= -1403673233;
assign addr[20748]= -1460659832;
assign addr[20749]= -1515793473;
assign addr[20750]= -1569004214;
assign addr[20751]= -1620224553;
assign addr[20752]= -1669389513;
assign addr[20753]= -1716436725;
assign addr[20754]= -1761306505;
assign addr[20755]= -1803941934;
assign addr[20756]= -1844288924;
assign addr[20757]= -1882296293;
assign addr[20758]= -1917915825;
assign addr[20759]= -1951102334;
assign addr[20760]= -1981813720;
assign addr[20761]= -2010011024;
assign addr[20762]= -2035658475;
assign addr[20763]= -2058723538;
assign addr[20764]= -2079176953;
assign addr[20765]= -2096992772;
assign addr[20766]= -2112148396;
assign addr[20767]= -2124624598;
assign addr[20768]= -2134405552;
assign addr[20769]= -2141478848;
assign addr[20770]= -2145835515;
assign addr[20771]= -2147470025;
assign addr[20772]= -2146380306;
assign addr[20773]= -2142567738;
assign addr[20774]= -2136037160;
assign addr[20775]= -2126796855;
assign addr[20776]= -2114858546;
assign addr[20777]= -2100237377;
assign addr[20778]= -2082951896;
assign addr[20779]= -2063024031;
assign addr[20780]= -2040479063;
assign addr[20781]= -2015345591;
assign addr[20782]= -1987655498;
assign addr[20783]= -1957443913;
assign addr[20784]= -1924749160;
assign addr[20785]= -1889612716;
assign addr[20786]= -1852079154;
assign addr[20787]= -1812196087;
assign addr[20788]= -1770014111;
assign addr[20789]= -1725586737;
assign addr[20790]= -1678970324;
assign addr[20791]= -1630224009;
assign addr[20792]= -1579409630;
assign addr[20793]= -1526591649;
assign addr[20794]= -1471837070;
assign addr[20795]= -1415215352;
assign addr[20796]= -1356798326;
assign addr[20797]= -1296660098;
assign addr[20798]= -1234876957;
assign addr[20799]= -1171527280;
assign addr[20800]= -1106691431;
assign addr[20801]= -1040451659;
assign addr[20802]= -972891995;
assign addr[20803]= -904098143;
assign addr[20804]= -834157373;
assign addr[20805]= -763158411;
assign addr[20806]= -691191324;
assign addr[20807]= -618347408;
assign addr[20808]= -544719071;
assign addr[20809]= -470399716;
assign addr[20810]= -395483624;
assign addr[20811]= -320065829;
assign addr[20812]= -244242007;
assign addr[20813]= -168108346;
assign addr[20814]= -91761426;
assign addr[20815]= -15298099;
assign addr[20816]= 61184634;
assign addr[20817]= 137589750;
assign addr[20818]= 213820322;
assign addr[20819]= 289779648;
assign addr[20820]= 365371365;
assign addr[20821]= 440499581;
assign addr[20822]= 515068990;
assign addr[20823]= 588984994;
assign addr[20824]= 662153826;
assign addr[20825]= 734482665;
assign addr[20826]= 805879757;
assign addr[20827]= 876254528;
assign addr[20828]= 945517704;
assign addr[20829]= 1013581418;
assign addr[20830]= 1080359326;
assign addr[20831]= 1145766716;
assign addr[20832]= 1209720613;
assign addr[20833]= 1272139887;
assign addr[20834]= 1332945355;
assign addr[20835]= 1392059879;
assign addr[20836]= 1449408469;
assign addr[20837]= 1504918373;
assign addr[20838]= 1558519173;
assign addr[20839]= 1610142873;
assign addr[20840]= 1659723983;
assign addr[20841]= 1707199606;
assign addr[20842]= 1752509516;
assign addr[20843]= 1795596234;
assign addr[20844]= 1836405100;
assign addr[20845]= 1874884346;
assign addr[20846]= 1910985158;
assign addr[20847]= 1944661739;
assign addr[20848]= 1975871368;
assign addr[20849]= 2004574453;
assign addr[20850]= 2030734582;
assign addr[20851]= 2054318569;
assign addr[20852]= 2075296495;
assign addr[20853]= 2093641749;
assign addr[20854]= 2109331059;
assign addr[20855]= 2122344521;
assign addr[20856]= 2132665626;
assign addr[20857]= 2140281282;
assign addr[20858]= 2145181827;
assign addr[20859]= 2147361045;
assign addr[20860]= 2146816171;
assign addr[20861]= 2143547897;
assign addr[20862]= 2137560369;
assign addr[20863]= 2128861181;
assign addr[20864]= 2117461370;
assign addr[20865]= 2103375398;
assign addr[20866]= 2086621133;
assign addr[20867]= 2067219829;
assign addr[20868]= 2045196100;
assign addr[20869]= 2020577882;
assign addr[20870]= 1993396407;
assign addr[20871]= 1963686155;
assign addr[20872]= 1931484818;
assign addr[20873]= 1896833245;
assign addr[20874]= 1859775393;
assign addr[20875]= 1820358275;
assign addr[20876]= 1778631892;
assign addr[20877]= 1734649179;
assign addr[20878]= 1688465931;
assign addr[20879]= 1640140734;
assign addr[20880]= 1589734894;
assign addr[20881]= 1537312353;
assign addr[20882]= 1482939614;
assign addr[20883]= 1426685652;
assign addr[20884]= 1368621831;
assign addr[20885]= 1308821808;
assign addr[20886]= 1247361445;
assign addr[20887]= 1184318708;
assign addr[20888]= 1119773573;
assign addr[20889]= 1053807919;
assign addr[20890]= 986505429;
assign addr[20891]= 917951481;
assign addr[20892]= 848233042;
assign addr[20893]= 777438554;
assign addr[20894]= 705657826;
assign addr[20895]= 632981917;
assign addr[20896]= 559503022;
assign addr[20897]= 485314355;
assign addr[20898]= 410510029;
assign addr[20899]= 335184940;
assign addr[20900]= 259434643;
assign addr[20901]= 183355234;
assign addr[20902]= 107043224;
assign addr[20903]= 30595422;
assign addr[20904]= -45891193;
assign addr[20905]= -122319591;
assign addr[20906]= -198592817;
assign addr[20907]= -274614114;
assign addr[20908]= -350287041;
assign addr[20909]= -425515602;
assign addr[20910]= -500204365;
assign addr[20911]= -574258580;
assign addr[20912]= -647584304;
assign addr[20913]= -720088517;
assign addr[20914]= -791679244;
assign addr[20915]= -862265664;
assign addr[20916]= -931758235;
assign addr[20917]= -1000068799;
assign addr[20918]= -1067110699;
assign addr[20919]= -1132798888;
assign addr[20920]= -1197050035;
assign addr[20921]= -1259782632;
assign addr[20922]= -1320917099;
assign addr[20923]= -1380375881;
assign addr[20924]= -1438083551;
assign addr[20925]= -1493966902;
assign addr[20926]= -1547955041;
assign addr[20927]= -1599979481;
assign addr[20928]= -1649974225;
assign addr[20929]= -1697875851;
assign addr[20930]= -1743623590;
assign addr[20931]= -1787159411;
assign addr[20932]= -1828428082;
assign addr[20933]= -1867377253;
assign addr[20934]= -1903957513;
assign addr[20935]= -1938122457;
assign addr[20936]= -1969828744;
assign addr[20937]= -1999036154;
assign addr[20938]= -2025707632;
assign addr[20939]= -2049809346;
assign addr[20940]= -2071310720;
assign addr[20941]= -2090184478;
assign addr[20942]= -2106406677;
assign addr[20943]= -2119956737;
assign addr[20944]= -2130817471;
assign addr[20945]= -2138975100;
assign addr[20946]= -2144419275;
assign addr[20947]= -2147143090;
assign addr[20948]= -2147143090;
assign addr[20949]= -2144419275;
assign addr[20950]= -2138975100;
assign addr[20951]= -2130817471;
assign addr[20952]= -2119956737;
assign addr[20953]= -2106406677;
assign addr[20954]= -2090184478;
assign addr[20955]= -2071310720;
assign addr[20956]= -2049809346;
assign addr[20957]= -2025707632;
assign addr[20958]= -1999036154;
assign addr[20959]= -1969828744;
assign addr[20960]= -1938122457;
assign addr[20961]= -1903957513;
assign addr[20962]= -1867377253;
assign addr[20963]= -1828428082;
assign addr[20964]= -1787159411;
assign addr[20965]= -1743623590;
assign addr[20966]= -1697875851;
assign addr[20967]= -1649974225;
assign addr[20968]= -1599979481;
assign addr[20969]= -1547955041;
assign addr[20970]= -1493966902;
assign addr[20971]= -1438083551;
assign addr[20972]= -1380375881;
assign addr[20973]= -1320917099;
assign addr[20974]= -1259782632;
assign addr[20975]= -1197050035;
assign addr[20976]= -1132798888;
assign addr[20977]= -1067110699;
assign addr[20978]= -1000068799;
assign addr[20979]= -931758235;
assign addr[20980]= -862265664;
assign addr[20981]= -791679244;
assign addr[20982]= -720088517;
assign addr[20983]= -647584304;
assign addr[20984]= -574258580;
assign addr[20985]= -500204365;
assign addr[20986]= -425515602;
assign addr[20987]= -350287041;
assign addr[20988]= -274614114;
assign addr[20989]= -198592817;
assign addr[20990]= -122319591;
assign addr[20991]= -45891193;
assign addr[20992]= 30595422;
assign addr[20993]= 107043224;
assign addr[20994]= 183355234;
assign addr[20995]= 259434643;
assign addr[20996]= 335184940;
assign addr[20997]= 410510029;
assign addr[20998]= 485314355;
assign addr[20999]= 559503022;
assign addr[21000]= 632981917;
assign addr[21001]= 705657826;
assign addr[21002]= 777438554;
assign addr[21003]= 848233042;
assign addr[21004]= 917951481;
assign addr[21005]= 986505429;
assign addr[21006]= 1053807919;
assign addr[21007]= 1119773573;
assign addr[21008]= 1184318708;
assign addr[21009]= 1247361445;
assign addr[21010]= 1308821808;
assign addr[21011]= 1368621831;
assign addr[21012]= 1426685652;
assign addr[21013]= 1482939614;
assign addr[21014]= 1537312353;
assign addr[21015]= 1589734894;
assign addr[21016]= 1640140734;
assign addr[21017]= 1688465931;
assign addr[21018]= 1734649179;
assign addr[21019]= 1778631892;
assign addr[21020]= 1820358275;
assign addr[21021]= 1859775393;
assign addr[21022]= 1896833245;
assign addr[21023]= 1931484818;
assign addr[21024]= 1963686155;
assign addr[21025]= 1993396407;
assign addr[21026]= 2020577882;
assign addr[21027]= 2045196100;
assign addr[21028]= 2067219829;
assign addr[21029]= 2086621133;
assign addr[21030]= 2103375398;
assign addr[21031]= 2117461370;
assign addr[21032]= 2128861181;
assign addr[21033]= 2137560369;
assign addr[21034]= 2143547897;
assign addr[21035]= 2146816171;
assign addr[21036]= 2147361045;
assign addr[21037]= 2145181827;
assign addr[21038]= 2140281282;
assign addr[21039]= 2132665626;
assign addr[21040]= 2122344521;
assign addr[21041]= 2109331059;
assign addr[21042]= 2093641749;
assign addr[21043]= 2075296495;
assign addr[21044]= 2054318569;
assign addr[21045]= 2030734582;
assign addr[21046]= 2004574453;
assign addr[21047]= 1975871368;
assign addr[21048]= 1944661739;
assign addr[21049]= 1910985158;
assign addr[21050]= 1874884346;
assign addr[21051]= 1836405100;
assign addr[21052]= 1795596234;
assign addr[21053]= 1752509516;
assign addr[21054]= 1707199606;
assign addr[21055]= 1659723983;
assign addr[21056]= 1610142873;
assign addr[21057]= 1558519173;
assign addr[21058]= 1504918373;
assign addr[21059]= 1449408469;
assign addr[21060]= 1392059879;
assign addr[21061]= 1332945355;
assign addr[21062]= 1272139887;
assign addr[21063]= 1209720613;
assign addr[21064]= 1145766716;
assign addr[21065]= 1080359326;
assign addr[21066]= 1013581418;
assign addr[21067]= 945517704;
assign addr[21068]= 876254528;
assign addr[21069]= 805879757;
assign addr[21070]= 734482665;
assign addr[21071]= 662153826;
assign addr[21072]= 588984994;
assign addr[21073]= 515068990;
assign addr[21074]= 440499581;
assign addr[21075]= 365371365;
assign addr[21076]= 289779648;
assign addr[21077]= 213820322;
assign addr[21078]= 137589750;
assign addr[21079]= 61184634;
assign addr[21080]= -15298099;
assign addr[21081]= -91761426;
assign addr[21082]= -168108346;
assign addr[21083]= -244242007;
assign addr[21084]= -320065829;
assign addr[21085]= -395483624;
assign addr[21086]= -470399716;
assign addr[21087]= -544719071;
assign addr[21088]= -618347408;
assign addr[21089]= -691191324;
assign addr[21090]= -763158411;
assign addr[21091]= -834157373;
assign addr[21092]= -904098143;
assign addr[21093]= -972891995;
assign addr[21094]= -1040451659;
assign addr[21095]= -1106691431;
assign addr[21096]= -1171527280;
assign addr[21097]= -1234876957;
assign addr[21098]= -1296660098;
assign addr[21099]= -1356798326;
assign addr[21100]= -1415215352;
assign addr[21101]= -1471837070;
assign addr[21102]= -1526591649;
assign addr[21103]= -1579409630;
assign addr[21104]= -1630224009;
assign addr[21105]= -1678970324;
assign addr[21106]= -1725586737;
assign addr[21107]= -1770014111;
assign addr[21108]= -1812196087;
assign addr[21109]= -1852079154;
assign addr[21110]= -1889612716;
assign addr[21111]= -1924749160;
assign addr[21112]= -1957443913;
assign addr[21113]= -1987655498;
assign addr[21114]= -2015345591;
assign addr[21115]= -2040479063;
assign addr[21116]= -2063024031;
assign addr[21117]= -2082951896;
assign addr[21118]= -2100237377;
assign addr[21119]= -2114858546;
assign addr[21120]= -2126796855;
assign addr[21121]= -2136037160;
assign addr[21122]= -2142567738;
assign addr[21123]= -2146380306;
assign addr[21124]= -2147470025;
assign addr[21125]= -2145835515;
assign addr[21126]= -2141478848;
assign addr[21127]= -2134405552;
assign addr[21128]= -2124624598;
assign addr[21129]= -2112148396;
assign addr[21130]= -2096992772;
assign addr[21131]= -2079176953;
assign addr[21132]= -2058723538;
assign addr[21133]= -2035658475;
assign addr[21134]= -2010011024;
assign addr[21135]= -1981813720;
assign addr[21136]= -1951102334;
assign addr[21137]= -1917915825;
assign addr[21138]= -1882296293;
assign addr[21139]= -1844288924;
assign addr[21140]= -1803941934;
assign addr[21141]= -1761306505;
assign addr[21142]= -1716436725;
assign addr[21143]= -1669389513;
assign addr[21144]= -1620224553;
assign addr[21145]= -1569004214;
assign addr[21146]= -1515793473;
assign addr[21147]= -1460659832;
assign addr[21148]= -1403673233;
assign addr[21149]= -1344905966;
assign addr[21150]= -1284432584;
assign addr[21151]= -1222329801;
assign addr[21152]= -1158676398;
assign addr[21153]= -1093553126;
assign addr[21154]= -1027042599;
assign addr[21155]= -959229189;
assign addr[21156]= -890198924;
assign addr[21157]= -820039373;
assign addr[21158]= -748839539;
assign addr[21159]= -676689746;
assign addr[21160]= -603681519;
assign addr[21161]= -529907477;
assign addr[21162]= -455461206;
assign addr[21163]= -380437148;
assign addr[21164]= -304930476;
assign addr[21165]= -229036977;
assign addr[21166]= -152852926;
assign addr[21167]= -76474970;
assign addr[21168]= 0;
assign addr[21169]= 76474970;
assign addr[21170]= 152852926;
assign addr[21171]= 229036977;
assign addr[21172]= 304930476;
assign addr[21173]= 380437148;
assign addr[21174]= 455461206;
assign addr[21175]= 529907477;
assign addr[21176]= 603681519;
assign addr[21177]= 676689746;
assign addr[21178]= 748839539;
assign addr[21179]= 820039373;
assign addr[21180]= 890198924;
assign addr[21181]= 959229189;
assign addr[21182]= 1027042599;
assign addr[21183]= 1093553126;
assign addr[21184]= 1158676398;
assign addr[21185]= 1222329801;
assign addr[21186]= 1284432584;
assign addr[21187]= 1344905966;
assign addr[21188]= 1403673233;
assign addr[21189]= 1460659832;
assign addr[21190]= 1515793473;
assign addr[21191]= 1569004214;
assign addr[21192]= 1620224553;
assign addr[21193]= 1669389513;
assign addr[21194]= 1716436725;
assign addr[21195]= 1761306505;
assign addr[21196]= 1803941934;
assign addr[21197]= 1844288924;
assign addr[21198]= 1882296293;
assign addr[21199]= 1917915825;
assign addr[21200]= 1951102334;
assign addr[21201]= 1981813720;
assign addr[21202]= 2010011024;
assign addr[21203]= 2035658475;
assign addr[21204]= 2058723538;
assign addr[21205]= 2079176953;
assign addr[21206]= 2096992772;
assign addr[21207]= 2112148396;
assign addr[21208]= 2124624598;
assign addr[21209]= 2134405552;
assign addr[21210]= 2141478848;
assign addr[21211]= 2145835515;
assign addr[21212]= 2147470025;
assign addr[21213]= 2146380306;
assign addr[21214]= 2142567738;
assign addr[21215]= 2136037160;
assign addr[21216]= 2126796855;
assign addr[21217]= 2114858546;
assign addr[21218]= 2100237377;
assign addr[21219]= 2082951896;
assign addr[21220]= 2063024031;
assign addr[21221]= 2040479063;
assign addr[21222]= 2015345591;
assign addr[21223]= 1987655498;
assign addr[21224]= 1957443913;
assign addr[21225]= 1924749160;
assign addr[21226]= 1889612716;
assign addr[21227]= 1852079154;
assign addr[21228]= 1812196087;
assign addr[21229]= 1770014111;
assign addr[21230]= 1725586737;
assign addr[21231]= 1678970324;
assign addr[21232]= 1630224009;
assign addr[21233]= 1579409630;
assign addr[21234]= 1526591649;
assign addr[21235]= 1471837070;
assign addr[21236]= 1415215352;
assign addr[21237]= 1356798326;
assign addr[21238]= 1296660098;
assign addr[21239]= 1234876957;
assign addr[21240]= 1171527280;
assign addr[21241]= 1106691431;
assign addr[21242]= 1040451659;
assign addr[21243]= 972891995;
assign addr[21244]= 904098143;
assign addr[21245]= 834157373;
assign addr[21246]= 763158411;
assign addr[21247]= 691191324;
assign addr[21248]= 618347408;
assign addr[21249]= 544719071;
assign addr[21250]= 470399716;
assign addr[21251]= 395483624;
assign addr[21252]= 320065829;
assign addr[21253]= 244242007;
assign addr[21254]= 168108346;
assign addr[21255]= 91761426;
assign addr[21256]= 15298099;
assign addr[21257]= -61184634;
assign addr[21258]= -137589750;
assign addr[21259]= -213820322;
assign addr[21260]= -289779648;
assign addr[21261]= -365371365;
assign addr[21262]= -440499581;
assign addr[21263]= -515068990;
assign addr[21264]= -588984994;
assign addr[21265]= -662153826;
assign addr[21266]= -734482665;
assign addr[21267]= -805879757;
assign addr[21268]= -876254528;
assign addr[21269]= -945517704;
assign addr[21270]= -1013581418;
assign addr[21271]= -1080359326;
assign addr[21272]= -1145766716;
assign addr[21273]= -1209720613;
assign addr[21274]= -1272139887;
assign addr[21275]= -1332945355;
assign addr[21276]= -1392059879;
assign addr[21277]= -1449408469;
assign addr[21278]= -1504918373;
assign addr[21279]= -1558519173;
assign addr[21280]= -1610142873;
assign addr[21281]= -1659723983;
assign addr[21282]= -1707199606;
assign addr[21283]= -1752509516;
assign addr[21284]= -1795596234;
assign addr[21285]= -1836405100;
assign addr[21286]= -1874884346;
assign addr[21287]= -1910985158;
assign addr[21288]= -1944661739;
assign addr[21289]= -1975871368;
assign addr[21290]= -2004574453;
assign addr[21291]= -2030734582;
assign addr[21292]= -2054318569;
assign addr[21293]= -2075296495;
assign addr[21294]= -2093641749;
assign addr[21295]= -2109331059;
assign addr[21296]= -2122344521;
assign addr[21297]= -2132665626;
assign addr[21298]= -2140281282;
assign addr[21299]= -2145181827;
assign addr[21300]= -2147361045;
assign addr[21301]= -2146816171;
assign addr[21302]= -2143547897;
assign addr[21303]= -2137560369;
assign addr[21304]= -2128861181;
assign addr[21305]= -2117461370;
assign addr[21306]= -2103375398;
assign addr[21307]= -2086621133;
assign addr[21308]= -2067219829;
assign addr[21309]= -2045196100;
assign addr[21310]= -2020577882;
assign addr[21311]= -1993396407;
assign addr[21312]= -1963686155;
assign addr[21313]= -1931484818;
assign addr[21314]= -1896833245;
assign addr[21315]= -1859775393;
assign addr[21316]= -1820358275;
assign addr[21317]= -1778631892;
assign addr[21318]= -1734649179;
assign addr[21319]= -1688465931;
assign addr[21320]= -1640140734;
assign addr[21321]= -1589734894;
assign addr[21322]= -1537312353;
assign addr[21323]= -1482939614;
assign addr[21324]= -1426685652;
assign addr[21325]= -1368621831;
assign addr[21326]= -1308821808;
assign addr[21327]= -1247361445;
assign addr[21328]= -1184318708;
assign addr[21329]= -1119773573;
assign addr[21330]= -1053807919;
assign addr[21331]= -986505429;
assign addr[21332]= -917951481;
assign addr[21333]= -848233042;
assign addr[21334]= -777438554;
assign addr[21335]= -705657826;
assign addr[21336]= -632981917;
assign addr[21337]= -559503022;
assign addr[21338]= -485314355;
assign addr[21339]= -410510029;
assign addr[21340]= -335184940;
assign addr[21341]= -259434643;
assign addr[21342]= -183355234;
assign addr[21343]= -107043224;
assign addr[21344]= -30595422;
assign addr[21345]= 45891193;
assign addr[21346]= 122319591;
assign addr[21347]= 198592817;
assign addr[21348]= 274614114;
assign addr[21349]= 350287041;
assign addr[21350]= 425515602;
assign addr[21351]= 500204365;
assign addr[21352]= 574258580;
assign addr[21353]= 647584304;
assign addr[21354]= 720088517;
assign addr[21355]= 791679244;
assign addr[21356]= 862265664;
assign addr[21357]= 931758235;
assign addr[21358]= 1000068799;
assign addr[21359]= 1067110699;
assign addr[21360]= 1132798888;
assign addr[21361]= 1197050035;
assign addr[21362]= 1259782632;
assign addr[21363]= 1320917099;
assign addr[21364]= 1380375881;
assign addr[21365]= 1438083551;
assign addr[21366]= 1493966902;
assign addr[21367]= 1547955041;
assign addr[21368]= 1599979481;
assign addr[21369]= 1649974225;
assign addr[21370]= 1697875851;
assign addr[21371]= 1743623590;
assign addr[21372]= 1787159411;
assign addr[21373]= 1828428082;
assign addr[21374]= 1867377253;
assign addr[21375]= 1903957513;
assign addr[21376]= 1938122457;
assign addr[21377]= 1969828744;
assign addr[21378]= 1999036154;
assign addr[21379]= 2025707632;
assign addr[21380]= 2049809346;
assign addr[21381]= 2071310720;
assign addr[21382]= 2090184478;
assign addr[21383]= 2106406677;
assign addr[21384]= 2119956737;
assign addr[21385]= 2130817471;
assign addr[21386]= 2138975100;
assign addr[21387]= 2144419275;
assign addr[21388]= 2147143090;
assign addr[21389]= 2147143090;
assign addr[21390]= 2144419275;
assign addr[21391]= 2138975100;
assign addr[21392]= 2130817471;
assign addr[21393]= 2119956737;
assign addr[21394]= 2106406677;
assign addr[21395]= 2090184478;
assign addr[21396]= 2071310720;
assign addr[21397]= 2049809346;
assign addr[21398]= 2025707632;
assign addr[21399]= 1999036154;
assign addr[21400]= 1969828744;
assign addr[21401]= 1938122457;
assign addr[21402]= 1903957513;
assign addr[21403]= 1867377253;
assign addr[21404]= 1828428082;
assign addr[21405]= 1787159411;
assign addr[21406]= 1743623590;
assign addr[21407]= 1697875851;
assign addr[21408]= 1649974225;
assign addr[21409]= 1599979481;
assign addr[21410]= 1547955041;
assign addr[21411]= 1493966902;
assign addr[21412]= 1438083551;
assign addr[21413]= 1380375881;
assign addr[21414]= 1320917099;
assign addr[21415]= 1259782632;
assign addr[21416]= 1197050035;
assign addr[21417]= 1132798888;
assign addr[21418]= 1067110699;
assign addr[21419]= 1000068799;
assign addr[21420]= 931758235;
assign addr[21421]= 862265664;
assign addr[21422]= 791679244;
assign addr[21423]= 720088517;
assign addr[21424]= 647584304;
assign addr[21425]= 574258580;
assign addr[21426]= 500204365;
assign addr[21427]= 425515602;
assign addr[21428]= 350287041;
assign addr[21429]= 274614114;
assign addr[21430]= 198592817;
assign addr[21431]= 122319591;
assign addr[21432]= 45891193;
assign addr[21433]= -30595422;
assign addr[21434]= -107043224;
assign addr[21435]= -183355234;
assign addr[21436]= -259434643;
assign addr[21437]= -335184940;
assign addr[21438]= -410510029;
assign addr[21439]= -485314355;
assign addr[21440]= -559503022;
assign addr[21441]= -632981917;
assign addr[21442]= -705657826;
assign addr[21443]= -777438554;
assign addr[21444]= -848233042;
assign addr[21445]= -917951481;
assign addr[21446]= -986505429;
assign addr[21447]= -1053807919;
assign addr[21448]= -1119773573;
assign addr[21449]= -1184318708;
assign addr[21450]= -1247361445;
assign addr[21451]= -1308821808;
assign addr[21452]= -1368621831;
assign addr[21453]= -1426685652;
assign addr[21454]= -1482939614;
assign addr[21455]= -1537312353;
assign addr[21456]= -1589734894;
assign addr[21457]= -1640140734;
assign addr[21458]= -1688465931;
assign addr[21459]= -1734649179;
assign addr[21460]= -1778631892;
assign addr[21461]= -1820358275;
assign addr[21462]= -1859775393;
assign addr[21463]= -1896833245;
assign addr[21464]= -1931484818;
assign addr[21465]= -1963686155;
assign addr[21466]= -1993396407;
assign addr[21467]= -2020577882;
assign addr[21468]= -2045196100;
assign addr[21469]= -2067219829;
assign addr[21470]= -2086621133;
assign addr[21471]= -2103375398;
assign addr[21472]= -2117461370;
assign addr[21473]= -2128861181;
assign addr[21474]= -2137560369;
assign addr[21475]= -2143547897;
assign addr[21476]= -2146816171;
assign addr[21477]= -2147361045;
assign addr[21478]= -2145181827;
assign addr[21479]= -2140281282;
assign addr[21480]= -2132665626;
assign addr[21481]= -2122344521;
assign addr[21482]= -2109331059;
assign addr[21483]= -2093641749;
assign addr[21484]= -2075296495;
assign addr[21485]= -2054318569;
assign addr[21486]= -2030734582;
assign addr[21487]= -2004574453;
assign addr[21488]= -1975871368;
assign addr[21489]= -1944661739;
assign addr[21490]= -1910985158;
assign addr[21491]= -1874884346;
assign addr[21492]= -1836405100;
assign addr[21493]= -1795596234;
assign addr[21494]= -1752509516;
assign addr[21495]= -1707199606;
assign addr[21496]= -1659723983;
assign addr[21497]= -1610142873;
assign addr[21498]= -1558519173;
assign addr[21499]= -1504918373;
assign addr[21500]= -1449408469;
assign addr[21501]= -1392059879;
assign addr[21502]= -1332945355;
assign addr[21503]= -1272139887;
assign addr[21504]= -1209720613;
assign addr[21505]= -1145766716;
assign addr[21506]= -1080359326;
assign addr[21507]= -1013581418;
assign addr[21508]= -945517704;
assign addr[21509]= -876254528;
assign addr[21510]= -805879757;
assign addr[21511]= -734482665;
assign addr[21512]= -662153826;
assign addr[21513]= -588984994;
assign addr[21514]= -515068990;
assign addr[21515]= -440499581;
assign addr[21516]= -365371365;
assign addr[21517]= -289779648;
assign addr[21518]= -213820322;
assign addr[21519]= -137589750;
assign addr[21520]= -61184634;
assign addr[21521]= 15298099;
assign addr[21522]= 91761426;
assign addr[21523]= 168108346;
assign addr[21524]= 244242007;
assign addr[21525]= 320065829;
assign addr[21526]= 395483624;
assign addr[21527]= 470399716;
assign addr[21528]= 544719071;
assign addr[21529]= 618347408;
assign addr[21530]= 691191324;
assign addr[21531]= 763158411;
assign addr[21532]= 834157373;
assign addr[21533]= 904098143;
assign addr[21534]= 972891995;
assign addr[21535]= 1040451659;
assign addr[21536]= 1106691431;
assign addr[21537]= 1171527280;
assign addr[21538]= 1234876957;
assign addr[21539]= 1296660098;
assign addr[21540]= 1356798326;
assign addr[21541]= 1415215352;
assign addr[21542]= 1471837070;
assign addr[21543]= 1526591649;
assign addr[21544]= 1579409630;
assign addr[21545]= 1630224009;
assign addr[21546]= 1678970324;
assign addr[21547]= 1725586737;
assign addr[21548]= 1770014111;
assign addr[21549]= 1812196087;
assign addr[21550]= 1852079154;
assign addr[21551]= 1889612716;
assign addr[21552]= 1924749160;
assign addr[21553]= 1957443913;
assign addr[21554]= 1987655498;
assign addr[21555]= 2015345591;
assign addr[21556]= 2040479063;
assign addr[21557]= 2063024031;
assign addr[21558]= 2082951896;
assign addr[21559]= 2100237377;
assign addr[21560]= 2114858546;
assign addr[21561]= 2126796855;
assign addr[21562]= 2136037160;
assign addr[21563]= 2142567738;
assign addr[21564]= 2146380306;
assign addr[21565]= 2147470025;
assign addr[21566]= 2145835515;
assign addr[21567]= 2141478848;
assign addr[21568]= 2134405552;
assign addr[21569]= 2124624598;
assign addr[21570]= 2112148396;
assign addr[21571]= 2096992772;
assign addr[21572]= 2079176953;
assign addr[21573]= 2058723538;
assign addr[21574]= 2035658475;
assign addr[21575]= 2010011024;
assign addr[21576]= 1981813720;
assign addr[21577]= 1951102334;
assign addr[21578]= 1917915825;
assign addr[21579]= 1882296293;
assign addr[21580]= 1844288924;
assign addr[21581]= 1803941934;
assign addr[21582]= 1761306505;
assign addr[21583]= 1716436725;
assign addr[21584]= 1669389513;
assign addr[21585]= 1620224553;
assign addr[21586]= 1569004214;
assign addr[21587]= 1515793473;
assign addr[21588]= 1460659832;
assign addr[21589]= 1403673233;
assign addr[21590]= 1344905966;
assign addr[21591]= 1284432584;
assign addr[21592]= 1222329801;
assign addr[21593]= 1158676398;
assign addr[21594]= 1093553126;
assign addr[21595]= 1027042599;
assign addr[21596]= 959229189;
assign addr[21597]= 890198924;
assign addr[21598]= 820039373;
assign addr[21599]= 748839539;
assign addr[21600]= 676689746;
assign addr[21601]= 603681519;
assign addr[21602]= 529907477;
assign addr[21603]= 455461206;
assign addr[21604]= 380437148;
assign addr[21605]= 304930476;
assign addr[21606]= 229036977;
assign addr[21607]= 152852926;
assign addr[21608]= 76474970;
assign addr[21609]= 0;
assign addr[21610]= -76474970;
assign addr[21611]= -152852926;
assign addr[21612]= -229036977;
assign addr[21613]= -304930476;
assign addr[21614]= -380437148;
assign addr[21615]= -455461206;
assign addr[21616]= -529907477;
assign addr[21617]= -603681519;
assign addr[21618]= -676689746;
assign addr[21619]= -748839539;
assign addr[21620]= -820039373;
assign addr[21621]= -890198924;
assign addr[21622]= -959229189;
assign addr[21623]= -1027042599;
assign addr[21624]= -1093553126;
assign addr[21625]= -1158676398;
assign addr[21626]= -1222329801;
assign addr[21627]= -1284432584;
assign addr[21628]= -1344905966;
assign addr[21629]= -1403673233;
assign addr[21630]= -1460659832;
assign addr[21631]= -1515793473;
assign addr[21632]= -1569004214;
assign addr[21633]= -1620224553;
assign addr[21634]= -1669389513;
assign addr[21635]= -1716436725;
assign addr[21636]= -1761306505;
assign addr[21637]= -1803941934;
assign addr[21638]= -1844288924;
assign addr[21639]= -1882296293;
assign addr[21640]= -1917915825;
assign addr[21641]= -1951102334;
assign addr[21642]= -1981813720;
assign addr[21643]= -2010011024;
assign addr[21644]= -2035658475;
assign addr[21645]= -2058723538;
assign addr[21646]= -2079176953;
assign addr[21647]= -2096992772;
assign addr[21648]= -2112148396;
assign addr[21649]= -2124624598;
assign addr[21650]= -2134405552;
assign addr[21651]= -2141478848;
assign addr[21652]= -2145835515;
assign addr[21653]= -2147470025;
assign addr[21654]= -2146380306;
assign addr[21655]= -2142567738;
assign addr[21656]= -2136037160;
assign addr[21657]= -2126796855;
assign addr[21658]= -2114858546;
assign addr[21659]= -2100237377;
assign addr[21660]= -2082951896;
assign addr[21661]= -2063024031;
assign addr[21662]= -2040479063;
assign addr[21663]= -2015345591;
assign addr[21664]= -1987655498;
assign addr[21665]= -1957443913;
assign addr[21666]= -1924749160;
assign addr[21667]= -1889612716;
assign addr[21668]= -1852079154;
assign addr[21669]= -1812196087;
assign addr[21670]= -1770014111;
assign addr[21671]= -1725586737;
assign addr[21672]= -1678970324;
assign addr[21673]= -1630224009;
assign addr[21674]= -1579409630;
assign addr[21675]= -1526591649;
assign addr[21676]= -1471837070;
assign addr[21677]= -1415215352;
assign addr[21678]= -1356798326;
assign addr[21679]= -1296660098;
assign addr[21680]= -1234876957;
assign addr[21681]= -1171527280;
assign addr[21682]= -1106691431;
assign addr[21683]= -1040451659;
assign addr[21684]= -972891995;
assign addr[21685]= -904098143;
assign addr[21686]= -834157373;
assign addr[21687]= -763158411;
assign addr[21688]= -691191324;
assign addr[21689]= -618347408;
assign addr[21690]= -544719071;
assign addr[21691]= -470399716;
assign addr[21692]= -395483624;
assign addr[21693]= -320065829;
assign addr[21694]= -244242007;
assign addr[21695]= -168108346;
assign addr[21696]= -91761426;
assign addr[21697]= -15298099;
assign addr[21698]= 61184634;
assign addr[21699]= 137589750;
assign addr[21700]= 213820322;
assign addr[21701]= 289779648;
assign addr[21702]= 365371365;
assign addr[21703]= 440499581;
assign addr[21704]= 515068990;
assign addr[21705]= 588984994;
assign addr[21706]= 662153826;
assign addr[21707]= 734482665;
assign addr[21708]= 805879757;
assign addr[21709]= 876254528;
assign addr[21710]= 945517704;
assign addr[21711]= 1013581418;
assign addr[21712]= 1080359326;
assign addr[21713]= 1145766716;
assign addr[21714]= 1209720613;
assign addr[21715]= 1272139887;
assign addr[21716]= 1332945355;
assign addr[21717]= 1392059879;
assign addr[21718]= 1449408469;
assign addr[21719]= 1504918373;
assign addr[21720]= 1558519173;
assign addr[21721]= 1610142873;
assign addr[21722]= 1659723983;
assign addr[21723]= 1707199606;
assign addr[21724]= 1752509516;
assign addr[21725]= 1795596234;
assign addr[21726]= 1836405100;
assign addr[21727]= 1874884346;
assign addr[21728]= 1910985158;
assign addr[21729]= 1944661739;
assign addr[21730]= 1975871368;
assign addr[21731]= 2004574453;
assign addr[21732]= 2030734582;
assign addr[21733]= 2054318569;
assign addr[21734]= 2075296495;
assign addr[21735]= 2093641749;
assign addr[21736]= 2109331059;
assign addr[21737]= 2122344521;
assign addr[21738]= 2132665626;
assign addr[21739]= 2140281282;
assign addr[21740]= 2145181827;
assign addr[21741]= 2147361045;
assign addr[21742]= 2146816171;
assign addr[21743]= 2143547897;
assign addr[21744]= 2137560369;
assign addr[21745]= 2128861181;
assign addr[21746]= 2117461370;
assign addr[21747]= 2103375398;
assign addr[21748]= 2086621133;
assign addr[21749]= 2067219829;
assign addr[21750]= 2045196100;
assign addr[21751]= 2020577882;
assign addr[21752]= 1993396407;
assign addr[21753]= 1963686155;
assign addr[21754]= 1931484818;
assign addr[21755]= 1896833245;
assign addr[21756]= 1859775393;
assign addr[21757]= 1820358275;
assign addr[21758]= 1778631892;
assign addr[21759]= 1734649179;
assign addr[21760]= 1688465931;
assign addr[21761]= 1640140734;
assign addr[21762]= 1589734894;
assign addr[21763]= 1537312353;
assign addr[21764]= 1482939614;
assign addr[21765]= 1426685652;
assign addr[21766]= 1368621831;
assign addr[21767]= 1308821808;
assign addr[21768]= 1247361445;
assign addr[21769]= 1184318708;
assign addr[21770]= 1119773573;
assign addr[21771]= 1053807919;
assign addr[21772]= 986505429;
assign addr[21773]= 917951481;
assign addr[21774]= 848233042;
assign addr[21775]= 777438554;
assign addr[21776]= 705657826;
assign addr[21777]= 632981917;
assign addr[21778]= 559503022;
assign addr[21779]= 485314355;
assign addr[21780]= 410510029;
assign addr[21781]= 335184940;
assign addr[21782]= 259434643;
assign addr[21783]= 183355234;
assign addr[21784]= 107043224;
assign addr[21785]= 30595422;
assign addr[21786]= -45891193;
assign addr[21787]= -122319591;
assign addr[21788]= -198592817;
assign addr[21789]= -274614114;
assign addr[21790]= -350287041;
assign addr[21791]= -425515602;
assign addr[21792]= -500204365;
assign addr[21793]= -574258580;
assign addr[21794]= -647584304;
assign addr[21795]= -720088517;
assign addr[21796]= -791679244;
assign addr[21797]= -862265664;
assign addr[21798]= -931758235;
assign addr[21799]= -1000068799;
assign addr[21800]= -1067110699;
assign addr[21801]= -1132798888;
assign addr[21802]= -1197050035;
assign addr[21803]= -1259782632;
assign addr[21804]= -1320917099;
assign addr[21805]= -1380375881;
assign addr[21806]= -1438083551;
assign addr[21807]= -1493966902;
assign addr[21808]= -1547955041;
assign addr[21809]= -1599979481;
assign addr[21810]= -1649974225;
assign addr[21811]= -1697875851;
assign addr[21812]= -1743623590;
assign addr[21813]= -1787159411;
assign addr[21814]= -1828428082;
assign addr[21815]= -1867377253;
assign addr[21816]= -1903957513;
assign addr[21817]= -1938122457;
assign addr[21818]= -1969828744;
assign addr[21819]= -1999036154;
assign addr[21820]= -2025707632;
assign addr[21821]= -2049809346;
assign addr[21822]= -2071310720;
assign addr[21823]= -2090184478;
assign addr[21824]= -2106406677;
assign addr[21825]= -2119956737;
assign addr[21826]= -2130817471;
assign addr[21827]= -2138975100;
assign addr[21828]= -2144419275;
assign addr[21829]= -2147143090;
assign addr[21830]= -2147143090;
assign addr[21831]= -2144419275;
assign addr[21832]= -2138975100;
assign addr[21833]= -2130817471;
assign addr[21834]= -2119956737;
assign addr[21835]= -2106406677;
assign addr[21836]= -2090184478;
assign addr[21837]= -2071310720;
assign addr[21838]= -2049809346;
assign addr[21839]= -2025707632;
assign addr[21840]= -1999036154;
assign addr[21841]= -1969828744;
assign addr[21842]= -1938122457;
assign addr[21843]= -1903957513;
assign addr[21844]= -1867377253;
assign addr[21845]= -1828428082;
assign addr[21846]= -1787159411;
assign addr[21847]= -1743623590;
assign addr[21848]= -1697875851;
assign addr[21849]= -1649974225;
assign addr[21850]= -1599979481;
assign addr[21851]= -1547955041;
assign addr[21852]= -1493966902;
assign addr[21853]= -1438083551;
assign addr[21854]= -1380375881;
assign addr[21855]= -1320917099;
assign addr[21856]= -1259782632;
assign addr[21857]= -1197050035;
assign addr[21858]= -1132798888;
assign addr[21859]= -1067110699;
assign addr[21860]= -1000068799;
assign addr[21861]= -931758235;
assign addr[21862]= -862265664;
assign addr[21863]= -791679244;
assign addr[21864]= -720088517;
assign addr[21865]= -647584304;
assign addr[21866]= -574258580;
assign addr[21867]= -500204365;
assign addr[21868]= -425515602;
assign addr[21869]= -350287041;
assign addr[21870]= -274614114;
assign addr[21871]= -198592817;
assign addr[21872]= -122319591;
assign addr[21873]= -45891193;
assign addr[21874]= 30595422;
assign addr[21875]= 107043224;
assign addr[21876]= 183355234;
assign addr[21877]= 259434643;
assign addr[21878]= 335184940;
assign addr[21879]= 410510029;
assign addr[21880]= 485314355;
assign addr[21881]= 559503022;
assign addr[21882]= 632981917;
assign addr[21883]= 705657826;
assign addr[21884]= 777438554;
assign addr[21885]= 848233042;
assign addr[21886]= 917951481;
assign addr[21887]= 986505429;
assign addr[21888]= 1053807919;
assign addr[21889]= 1119773573;
assign addr[21890]= 1184318708;
assign addr[21891]= 1247361445;
assign addr[21892]= 1308821808;
assign addr[21893]= 1368621831;
assign addr[21894]= 1426685652;
assign addr[21895]= 1482939614;
assign addr[21896]= 1537312353;
assign addr[21897]= 1589734894;
assign addr[21898]= 1640140734;
assign addr[21899]= 1688465931;
assign addr[21900]= 1734649179;
assign addr[21901]= 1778631892;
assign addr[21902]= 1820358275;
assign addr[21903]= 1859775393;
assign addr[21904]= 1896833245;
assign addr[21905]= 1931484818;
assign addr[21906]= 1963686155;
assign addr[21907]= 1993396407;
assign addr[21908]= 2020577882;
assign addr[21909]= 2045196100;
assign addr[21910]= 2067219829;
assign addr[21911]= 2086621133;
assign addr[21912]= 2103375398;
assign addr[21913]= 2117461370;
assign addr[21914]= 2128861181;
assign addr[21915]= 2137560369;
assign addr[21916]= 2143547897;
assign addr[21917]= 2146816171;
assign addr[21918]= 2147361045;
assign addr[21919]= 2145181827;
assign addr[21920]= 2140281282;
assign addr[21921]= 2132665626;
assign addr[21922]= 2122344521;
assign addr[21923]= 2109331059;
assign addr[21924]= 2093641749;
assign addr[21925]= 2075296495;
assign addr[21926]= 2054318569;
assign addr[21927]= 2030734582;
assign addr[21928]= 2004574453;
assign addr[21929]= 1975871368;
assign addr[21930]= 1944661739;
assign addr[21931]= 1910985158;
assign addr[21932]= 1874884346;
assign addr[21933]= 1836405100;
assign addr[21934]= 1795596234;
assign addr[21935]= 1752509516;
assign addr[21936]= 1707199606;
assign addr[21937]= 1659723983;
assign addr[21938]= 1610142873;
assign addr[21939]= 1558519173;
assign addr[21940]= 1504918373;
assign addr[21941]= 1449408469;
assign addr[21942]= 1392059879;
assign addr[21943]= 1332945355;
assign addr[21944]= 1272139887;
assign addr[21945]= 1209720613;
assign addr[21946]= 1145766716;
assign addr[21947]= 1080359326;
assign addr[21948]= 1013581418;
assign addr[21949]= 945517704;
assign addr[21950]= 876254528;
assign addr[21951]= 805879757;
assign addr[21952]= 734482665;
assign addr[21953]= 662153826;
assign addr[21954]= 588984994;
assign addr[21955]= 515068990;
assign addr[21956]= 440499581;
assign addr[21957]= 365371365;
assign addr[21958]= 289779648;
assign addr[21959]= 213820322;
assign addr[21960]= 137589750;
assign addr[21961]= 61184634;
assign addr[21962]= -15298099;
assign addr[21963]= -91761426;
assign addr[21964]= -168108346;
assign addr[21965]= -244242007;
assign addr[21966]= -320065829;
assign addr[21967]= -395483624;
assign addr[21968]= -470399716;
assign addr[21969]= -544719071;
assign addr[21970]= -618347408;
assign addr[21971]= -691191324;
assign addr[21972]= -763158411;
assign addr[21973]= -834157373;
assign addr[21974]= -904098143;
assign addr[21975]= -972891995;
assign addr[21976]= -1040451659;
assign addr[21977]= -1106691431;
assign addr[21978]= -1171527280;
assign addr[21979]= -1234876957;
assign addr[21980]= -1296660098;
assign addr[21981]= -1356798326;
assign addr[21982]= -1415215352;
assign addr[21983]= -1471837070;
assign addr[21984]= -1526591649;
assign addr[21985]= -1579409630;
assign addr[21986]= -1630224009;
assign addr[21987]= -1678970324;
assign addr[21988]= -1725586737;
assign addr[21989]= -1770014111;
assign addr[21990]= -1812196087;
assign addr[21991]= -1852079154;
assign addr[21992]= -1889612716;
assign addr[21993]= -1924749160;
assign addr[21994]= -1957443913;
assign addr[21995]= -1987655498;
assign addr[21996]= -2015345591;
assign addr[21997]= -2040479063;
assign addr[21998]= -2063024031;
assign addr[21999]= -2082951896;
assign addr[22000]= -2100237377;
assign addr[22001]= -2114858546;
assign addr[22002]= -2126796855;
assign addr[22003]= -2136037160;
assign addr[22004]= -2142567738;
assign addr[22005]= -2146380306;
assign addr[22006]= -2147470025;
assign addr[22007]= -2145835515;
assign addr[22008]= -2141478848;
assign addr[22009]= -2134405552;
assign addr[22010]= -2124624598;
assign addr[22011]= -2112148396;
assign addr[22012]= -2096992772;
assign addr[22013]= -2079176953;
assign addr[22014]= -2058723538;
assign addr[22015]= -2035658475;
assign addr[22016]= -2010011024;
assign addr[22017]= -1981813720;
assign addr[22018]= -1951102334;
assign addr[22019]= -1917915825;
assign addr[22020]= -1882296293;
assign addr[22021]= -1844288924;
assign addr[22022]= -1803941934;
assign addr[22023]= -1761306505;
assign addr[22024]= -1716436725;
assign addr[22025]= -1669389513;
assign addr[22026]= -1620224553;
assign addr[22027]= -1569004214;
assign addr[22028]= -1515793473;
assign addr[22029]= -1460659832;
assign addr[22030]= -1403673233;
assign addr[22031]= -1344905966;
assign addr[22032]= -1284432584;
assign addr[22033]= -1222329801;
assign addr[22034]= -1158676398;
assign addr[22035]= -1093553126;
assign addr[22036]= -1027042599;
assign addr[22037]= -959229189;
assign addr[22038]= -890198924;
assign addr[22039]= -820039373;
assign addr[22040]= -748839539;
assign addr[22041]= -676689746;
assign addr[22042]= -603681519;
assign addr[22043]= -529907477;
assign addr[22044]= -455461206;
assign addr[22045]= -380437148;
assign addr[22046]= -304930476;
assign addr[22047]= -229036977;
assign addr[22048]= -152852926;
assign addr[22049]= -76474970;
assign addr[22050]= 0;
assign addr[22051]= 76474970;
assign addr[22052]= 152852926;
assign addr[22053]= 229036977;
assign addr[22054]= 304930476;
assign addr[22055]= 380437148;
assign addr[22056]= 455461206;
assign addr[22057]= 529907477;
assign addr[22058]= 603681519;
assign addr[22059]= 676689746;
assign addr[22060]= 748839539;
assign addr[22061]= 820039373;
assign addr[22062]= 890198924;
assign addr[22063]= 959229189;
assign addr[22064]= 1027042599;
assign addr[22065]= 1093553126;
assign addr[22066]= 1158676398;
assign addr[22067]= 1222329801;
assign addr[22068]= 1284432584;
assign addr[22069]= 1344905966;
assign addr[22070]= 1403673233;
assign addr[22071]= 1460659832;
assign addr[22072]= 1515793473;
assign addr[22073]= 1569004214;
assign addr[22074]= 1620224553;
assign addr[22075]= 1669389513;
assign addr[22076]= 1716436725;
assign addr[22077]= 1761306505;
assign addr[22078]= 1803941934;
assign addr[22079]= 1844288924;
assign addr[22080]= 1882296293;
assign addr[22081]= 1917915825;
assign addr[22082]= 1951102334;
assign addr[22083]= 1981813720;
assign addr[22084]= 2010011024;
assign addr[22085]= 2035658475;
assign addr[22086]= 2058723538;
assign addr[22087]= 2079176953;
assign addr[22088]= 2096992772;
assign addr[22089]= 2112148396;
assign addr[22090]= 2124624598;
assign addr[22091]= 2134405552;
assign addr[22092]= 2141478848;
assign addr[22093]= 2145835515;
assign addr[22094]= 2147470025;
assign addr[22095]= 2146380306;
assign addr[22096]= 2142567738;
assign addr[22097]= 2136037160;
assign addr[22098]= 2126796855;
assign addr[22099]= 2114858546;
assign addr[22100]= 2100237377;
assign addr[22101]= 2082951896;
assign addr[22102]= 2063024031;
assign addr[22103]= 2040479063;
assign addr[22104]= 2015345591;
assign addr[22105]= 1987655498;
assign addr[22106]= 1957443913;
assign addr[22107]= 1924749160;
assign addr[22108]= 1889612716;
assign addr[22109]= 1852079154;
assign addr[22110]= 1812196087;
assign addr[22111]= 1770014111;
assign addr[22112]= 1725586737;
assign addr[22113]= 1678970324;
assign addr[22114]= 1630224009;
assign addr[22115]= 1579409630;
assign addr[22116]= 1526591649;
assign addr[22117]= 1471837070;
assign addr[22118]= 1415215352;
assign addr[22119]= 1356798326;
assign addr[22120]= 1296660098;
assign addr[22121]= 1234876957;
assign addr[22122]= 1171527280;
assign addr[22123]= 1106691431;
assign addr[22124]= 1040451659;
assign addr[22125]= 972891995;
assign addr[22126]= 904098143;
assign addr[22127]= 834157373;
assign addr[22128]= 763158411;
assign addr[22129]= 691191324;
assign addr[22130]= 618347408;
assign addr[22131]= 544719071;
assign addr[22132]= 470399716;
assign addr[22133]= 395483624;
assign addr[22134]= 320065829;
assign addr[22135]= 244242007;
assign addr[22136]= 168108346;
assign addr[22137]= 91761426;
assign addr[22138]= 15298099;
assign addr[22139]= -61184634;
assign addr[22140]= -137589750;
assign addr[22141]= -213820322;
assign addr[22142]= -289779648;
assign addr[22143]= -365371365;
assign addr[22144]= -440499581;
assign addr[22145]= -515068990;
assign addr[22146]= -588984994;
assign addr[22147]= -662153826;
assign addr[22148]= -734482665;
assign addr[22149]= -805879757;
assign addr[22150]= -876254528;
assign addr[22151]= -945517704;
assign addr[22152]= -1013581418;
assign addr[22153]= -1080359326;
assign addr[22154]= -1145766716;
assign addr[22155]= -1209720613;
assign addr[22156]= -1272139887;
assign addr[22157]= -1332945355;
assign addr[22158]= -1392059879;
assign addr[22159]= -1449408469;
assign addr[22160]= -1504918373;
assign addr[22161]= -1558519173;
assign addr[22162]= -1610142873;
assign addr[22163]= -1659723983;
assign addr[22164]= -1707199606;
assign addr[22165]= -1752509516;
assign addr[22166]= -1795596234;
assign addr[22167]= -1836405100;
assign addr[22168]= -1874884346;
assign addr[22169]= -1910985158;
assign addr[22170]= -1944661739;
assign addr[22171]= -1975871368;
assign addr[22172]= -2004574453;
assign addr[22173]= -2030734582;
assign addr[22174]= -2054318569;
assign addr[22175]= -2075296495;
assign addr[22176]= -2093641749;
assign addr[22177]= -2109331059;
assign addr[22178]= -2122344521;
assign addr[22179]= -2132665626;
assign addr[22180]= -2140281282;
assign addr[22181]= -2145181827;
assign addr[22182]= -2147361045;
assign addr[22183]= -2146816171;
assign addr[22184]= -2143547897;
assign addr[22185]= -2137560369;
assign addr[22186]= -2128861181;
assign addr[22187]= -2117461370;
assign addr[22188]= -2103375398;
assign addr[22189]= -2086621133;
assign addr[22190]= -2067219829;
assign addr[22191]= -2045196100;
assign addr[22192]= -2020577882;
assign addr[22193]= -1993396407;
assign addr[22194]= -1963686155;
assign addr[22195]= -1931484818;
assign addr[22196]= -1896833245;
assign addr[22197]= -1859775393;
assign addr[22198]= -1820358275;
assign addr[22199]= -1778631892;
assign addr[22200]= -1734649179;
assign addr[22201]= -1688465931;
assign addr[22202]= -1640140734;
assign addr[22203]= -1589734894;
assign addr[22204]= -1537312353;
assign addr[22205]= -1482939614;
assign addr[22206]= -1426685652;
assign addr[22207]= -1368621831;
assign addr[22208]= -1308821808;
assign addr[22209]= -1247361445;
assign addr[22210]= -1184318708;
assign addr[22211]= -1119773573;
assign addr[22212]= -1053807919;
assign addr[22213]= -986505429;
assign addr[22214]= -917951481;
assign addr[22215]= -848233042;
assign addr[22216]= -777438554;
assign addr[22217]= -705657826;
assign addr[22218]= -632981917;
assign addr[22219]= -559503022;
assign addr[22220]= -485314355;
assign addr[22221]= -410510029;
assign addr[22222]= -335184940;
assign addr[22223]= -259434643;
assign addr[22224]= -183355234;
assign addr[22225]= -107043224;
assign addr[22226]= -30595422;
assign addr[22227]= 45891193;
assign addr[22228]= 122319591;
assign addr[22229]= 198592817;
assign addr[22230]= 274614114;
assign addr[22231]= 350287041;
assign addr[22232]= 425515602;
assign addr[22233]= 500204365;
assign addr[22234]= 574258580;
assign addr[22235]= 647584304;
assign addr[22236]= 720088517;
assign addr[22237]= 791679244;
assign addr[22238]= 862265664;
assign addr[22239]= 931758235;
assign addr[22240]= 1000068799;
assign addr[22241]= 1067110699;
assign addr[22242]= 1132798888;
assign addr[22243]= 1197050035;
assign addr[22244]= 1259782632;
assign addr[22245]= 1320917099;
assign addr[22246]= 1380375881;
assign addr[22247]= 1438083551;
assign addr[22248]= 1493966902;
assign addr[22249]= 1547955041;
assign addr[22250]= 1599979481;
assign addr[22251]= 1649974225;
assign addr[22252]= 1697875851;
assign addr[22253]= 1743623590;
assign addr[22254]= 1787159411;
assign addr[22255]= 1828428082;
assign addr[22256]= 1867377253;
assign addr[22257]= 1903957513;
assign addr[22258]= 1938122457;
assign addr[22259]= 1969828744;
assign addr[22260]= 1999036154;
assign addr[22261]= 2025707632;
assign addr[22262]= 2049809346;
assign addr[22263]= 2071310720;
assign addr[22264]= 2090184478;
assign addr[22265]= 2106406677;
assign addr[22266]= 2119956737;
assign addr[22267]= 2130817471;
assign addr[22268]= 2138975100;
assign addr[22269]= 2144419275;
assign addr[22270]= 2147143090;
assign addr[22271]= 2147143090;
assign addr[22272]= 2144419275;
assign addr[22273]= 2138975100;
assign addr[22274]= 2130817471;
assign addr[22275]= 2119956737;
assign addr[22276]= 2106406677;
assign addr[22277]= 2090184478;
assign addr[22278]= 2071310720;
assign addr[22279]= 2049809346;
assign addr[22280]= 2025707632;
assign addr[22281]= 1999036154;
assign addr[22282]= 1969828744;
assign addr[22283]= 1938122457;
assign addr[22284]= 1903957513;
assign addr[22285]= 1867377253;
assign addr[22286]= 1828428082;
assign addr[22287]= 1787159411;
assign addr[22288]= 1743623590;
assign addr[22289]= 1697875851;
assign addr[22290]= 1649974225;
assign addr[22291]= 1599979481;
assign addr[22292]= 1547955041;
assign addr[22293]= 1493966902;
assign addr[22294]= 1438083551;
assign addr[22295]= 1380375881;
assign addr[22296]= 1320917099;
assign addr[22297]= 1259782632;
assign addr[22298]= 1197050035;
assign addr[22299]= 1132798888;
assign addr[22300]= 1067110699;
assign addr[22301]= 1000068799;
assign addr[22302]= 931758235;
assign addr[22303]= 862265664;
assign addr[22304]= 791679244;
assign addr[22305]= 720088517;
assign addr[22306]= 647584304;
assign addr[22307]= 574258580;
assign addr[22308]= 500204365;
assign addr[22309]= 425515602;
assign addr[22310]= 350287041;
assign addr[22311]= 274614114;
assign addr[22312]= 198592817;
assign addr[22313]= 122319591;
assign addr[22314]= 45891193;
assign addr[22315]= -30595422;
assign addr[22316]= -107043224;
assign addr[22317]= -183355234;
assign addr[22318]= -259434643;
assign addr[22319]= -335184940;
assign addr[22320]= -410510029;
assign addr[22321]= -485314355;
assign addr[22322]= -559503022;
assign addr[22323]= -632981917;
assign addr[22324]= -705657826;
assign addr[22325]= -777438554;
assign addr[22326]= -848233042;
assign addr[22327]= -917951481;
assign addr[22328]= -986505429;
assign addr[22329]= -1053807919;
assign addr[22330]= -1119773573;
assign addr[22331]= -1184318708;
assign addr[22332]= -1247361445;
assign addr[22333]= -1308821808;
assign addr[22334]= -1368621831;
assign addr[22335]= -1426685652;
assign addr[22336]= -1482939614;
assign addr[22337]= -1537312353;
assign addr[22338]= -1589734894;
assign addr[22339]= -1640140734;
assign addr[22340]= -1688465931;
assign addr[22341]= -1734649179;
assign addr[22342]= -1778631892;
assign addr[22343]= -1820358275;
assign addr[22344]= -1859775393;
assign addr[22345]= -1896833245;
assign addr[22346]= -1931484818;
assign addr[22347]= -1963686155;
assign addr[22348]= -1993396407;
assign addr[22349]= -2020577882;
assign addr[22350]= -2045196100;
assign addr[22351]= -2067219829;
assign addr[22352]= -2086621133;
assign addr[22353]= -2103375398;
assign addr[22354]= -2117461370;
assign addr[22355]= -2128861181;
assign addr[22356]= -2137560369;
assign addr[22357]= -2143547897;
assign addr[22358]= -2146816171;
assign addr[22359]= -2147361045;
assign addr[22360]= -2145181827;
assign addr[22361]= -2140281282;
assign addr[22362]= -2132665626;
assign addr[22363]= -2122344521;
assign addr[22364]= -2109331059;
assign addr[22365]= -2093641749;
assign addr[22366]= -2075296495;
assign addr[22367]= -2054318569;
assign addr[22368]= -2030734582;
assign addr[22369]= -2004574453;
assign addr[22370]= -1975871368;
assign addr[22371]= -1944661739;
assign addr[22372]= -1910985158;
assign addr[22373]= -1874884346;
assign addr[22374]= -1836405100;
assign addr[22375]= -1795596234;
assign addr[22376]= -1752509516;
assign addr[22377]= -1707199606;
assign addr[22378]= -1659723983;
assign addr[22379]= -1610142873;
assign addr[22380]= -1558519173;
assign addr[22381]= -1504918373;
assign addr[22382]= -1449408469;
assign addr[22383]= -1392059879;
assign addr[22384]= -1332945355;
assign addr[22385]= -1272139887;
assign addr[22386]= -1209720613;
assign addr[22387]= -1145766716;
assign addr[22388]= -1080359326;
assign addr[22389]= -1013581418;
assign addr[22390]= -945517704;
assign addr[22391]= -876254528;
assign addr[22392]= -805879757;
assign addr[22393]= -734482665;
assign addr[22394]= -662153826;
assign addr[22395]= -588984994;
assign addr[22396]= -515068990;
assign addr[22397]= -440499581;
assign addr[22398]= -365371365;
assign addr[22399]= -289779648;
assign addr[22400]= -213820322;
assign addr[22401]= -137589750;
assign addr[22402]= -61184634;
assign addr[22403]= 15298099;
assign addr[22404]= 91761426;
assign addr[22405]= 168108346;
assign addr[22406]= 244242007;
assign addr[22407]= 320065829;
assign addr[22408]= 395483624;
assign addr[22409]= 470399716;
assign addr[22410]= 544719071;
assign addr[22411]= 618347408;
assign addr[22412]= 691191324;
assign addr[22413]= 763158411;
assign addr[22414]= 834157373;
assign addr[22415]= 904098143;
assign addr[22416]= 972891995;
assign addr[22417]= 1040451659;
assign addr[22418]= 1106691431;
assign addr[22419]= 1171527280;
assign addr[22420]= 1234876957;
assign addr[22421]= 1296660098;
assign addr[22422]= 1356798326;
assign addr[22423]= 1415215352;
assign addr[22424]= 1471837070;
assign addr[22425]= 1526591649;
assign addr[22426]= 1579409630;
assign addr[22427]= 1630224009;
assign addr[22428]= 1678970324;
assign addr[22429]= 1725586737;
assign addr[22430]= 1770014111;
assign addr[22431]= 1812196087;
assign addr[22432]= 1852079154;
assign addr[22433]= 1889612716;
assign addr[22434]= 1924749160;
assign addr[22435]= 1957443913;
assign addr[22436]= 1987655498;
assign addr[22437]= 2015345591;
assign addr[22438]= 2040479063;
assign addr[22439]= 2063024031;
assign addr[22440]= 2082951896;
assign addr[22441]= 2100237377;
assign addr[22442]= 2114858546;
assign addr[22443]= 2126796855;
assign addr[22444]= 2136037160;
assign addr[22445]= 2142567738;
assign addr[22446]= 2146380306;
assign addr[22447]= 2147470025;
assign addr[22448]= 2145835515;
assign addr[22449]= 2141478848;
assign addr[22450]= 2134405552;
assign addr[22451]= 2124624598;
assign addr[22452]= 2112148396;
assign addr[22453]= 2096992772;
assign addr[22454]= 2079176953;
assign addr[22455]= 2058723538;
assign addr[22456]= 2035658475;
assign addr[22457]= 2010011024;
assign addr[22458]= 1981813720;
assign addr[22459]= 1951102334;
assign addr[22460]= 1917915825;
assign addr[22461]= 1882296293;
assign addr[22462]= 1844288924;
assign addr[22463]= 1803941934;
assign addr[22464]= 1761306505;
assign addr[22465]= 1716436725;
assign addr[22466]= 1669389513;
assign addr[22467]= 1620224553;
assign addr[22468]= 1569004214;
assign addr[22469]= 1515793473;
assign addr[22470]= 1460659832;
assign addr[22471]= 1403673233;
assign addr[22472]= 1344905966;
assign addr[22473]= 1284432584;
assign addr[22474]= 1222329801;
assign addr[22475]= 1158676398;
assign addr[22476]= 1093553126;
assign addr[22477]= 1027042599;
assign addr[22478]= 959229189;
assign addr[22479]= 890198924;
assign addr[22480]= 820039373;
assign addr[22481]= 748839539;
assign addr[22482]= 676689746;
assign addr[22483]= 603681519;
assign addr[22484]= 529907477;
assign addr[22485]= 455461206;
assign addr[22486]= 380437148;
assign addr[22487]= 304930476;
assign addr[22488]= 229036977;
assign addr[22489]= 152852926;
assign addr[22490]= 76474970;
assign addr[22491]= 0;
assign addr[22492]= -76474970;
assign addr[22493]= -152852926;
assign addr[22494]= -229036977;
assign addr[22495]= -304930476;
assign addr[22496]= -380437148;
assign addr[22497]= -455461206;
assign addr[22498]= -529907477;
assign addr[22499]= -603681519;
assign addr[22500]= -676689746;
assign addr[22501]= -748839539;
assign addr[22502]= -820039373;
assign addr[22503]= -890198924;
assign addr[22504]= -959229189;
assign addr[22505]= -1027042599;
assign addr[22506]= -1093553126;
assign addr[22507]= -1158676398;
assign addr[22508]= -1222329801;
assign addr[22509]= -1284432584;
assign addr[22510]= -1344905966;
assign addr[22511]= -1403673233;
assign addr[22512]= -1460659832;
assign addr[22513]= -1515793473;
assign addr[22514]= -1569004214;
assign addr[22515]= -1620224553;
assign addr[22516]= -1669389513;
assign addr[22517]= -1716436725;
assign addr[22518]= -1761306505;
assign addr[22519]= -1803941934;
assign addr[22520]= -1844288924;
assign addr[22521]= -1882296293;
assign addr[22522]= -1917915825;
assign addr[22523]= -1951102334;
assign addr[22524]= -1981813720;
assign addr[22525]= -2010011024;
assign addr[22526]= -2035658475;
assign addr[22527]= -2058723538;
assign addr[22528]= -2079176953;
assign addr[22529]= -2096992772;
assign addr[22530]= -2112148396;
assign addr[22531]= -2124624598;
assign addr[22532]= -2134405552;
assign addr[22533]= -2141478848;
assign addr[22534]= -2145835515;
assign addr[22535]= -2147470025;
assign addr[22536]= -2146380306;
assign addr[22537]= -2142567738;
assign addr[22538]= -2136037160;
assign addr[22539]= -2126796855;
assign addr[22540]= -2114858546;
assign addr[22541]= -2100237377;
assign addr[22542]= -2082951896;
assign addr[22543]= -2063024031;
assign addr[22544]= -2040479063;
assign addr[22545]= -2015345591;
assign addr[22546]= -1987655498;
assign addr[22547]= -1957443913;
assign addr[22548]= -1924749160;
assign addr[22549]= -1889612716;
assign addr[22550]= -1852079154;
assign addr[22551]= -1812196087;
assign addr[22552]= -1770014111;
assign addr[22553]= -1725586737;
assign addr[22554]= -1678970324;
assign addr[22555]= -1630224009;
assign addr[22556]= -1579409630;
assign addr[22557]= -1526591649;
assign addr[22558]= -1471837070;
assign addr[22559]= -1415215352;
assign addr[22560]= -1356798326;
assign addr[22561]= -1296660098;
assign addr[22562]= -1234876957;
assign addr[22563]= -1171527280;
assign addr[22564]= -1106691431;
assign addr[22565]= -1040451659;
assign addr[22566]= -972891995;
assign addr[22567]= -904098143;
assign addr[22568]= -834157373;
assign addr[22569]= -763158411;
assign addr[22570]= -691191324;
assign addr[22571]= -618347408;
assign addr[22572]= -544719071;
assign addr[22573]= -470399716;
assign addr[22574]= -395483624;
assign addr[22575]= -320065829;
assign addr[22576]= -244242007;
assign addr[22577]= -168108346;
assign addr[22578]= -91761426;
assign addr[22579]= -15298099;
assign addr[22580]= 61184634;
assign addr[22581]= 137589750;
assign addr[22582]= 213820322;
assign addr[22583]= 289779648;
assign addr[22584]= 365371365;
assign addr[22585]= 440499581;
assign addr[22586]= 515068990;
assign addr[22587]= 588984994;
assign addr[22588]= 662153826;
assign addr[22589]= 734482665;
assign addr[22590]= 805879757;
assign addr[22591]= 876254528;
assign addr[22592]= 945517704;
assign addr[22593]= 1013581418;
assign addr[22594]= 1080359326;
assign addr[22595]= 1145766716;
assign addr[22596]= 1209720613;
assign addr[22597]= 1272139887;
assign addr[22598]= 1332945355;
assign addr[22599]= 1392059879;
assign addr[22600]= 1449408469;
assign addr[22601]= 1504918373;
assign addr[22602]= 1558519173;
assign addr[22603]= 1610142873;
assign addr[22604]= 1659723983;
assign addr[22605]= 1707199606;
assign addr[22606]= 1752509516;
assign addr[22607]= 1795596234;
assign addr[22608]= 1836405100;
assign addr[22609]= 1874884346;
assign addr[22610]= 1910985158;
assign addr[22611]= 1944661739;
assign addr[22612]= 1975871368;
assign addr[22613]= 2004574453;
assign addr[22614]= 2030734582;
assign addr[22615]= 2054318569;
assign addr[22616]= 2075296495;
assign addr[22617]= 2093641749;
assign addr[22618]= 2109331059;
assign addr[22619]= 2122344521;
assign addr[22620]= 2132665626;
assign addr[22621]= 2140281282;
assign addr[22622]= 2145181827;
assign addr[22623]= 2147361045;
assign addr[22624]= 2146816171;
assign addr[22625]= 2143547897;
assign addr[22626]= 2137560369;
assign addr[22627]= 2128861181;
assign addr[22628]= 2117461370;
assign addr[22629]= 2103375398;
assign addr[22630]= 2086621133;
assign addr[22631]= 2067219829;
assign addr[22632]= 2045196100;
assign addr[22633]= 2020577882;
assign addr[22634]= 1993396407;
assign addr[22635]= 1963686155;
assign addr[22636]= 1931484818;
assign addr[22637]= 1896833245;
assign addr[22638]= 1859775393;
assign addr[22639]= 1820358275;
assign addr[22640]= 1778631892;
assign addr[22641]= 1734649179;
assign addr[22642]= 1688465931;
assign addr[22643]= 1640140734;
assign addr[22644]= 1589734894;
assign addr[22645]= 1537312353;
assign addr[22646]= 1482939614;
assign addr[22647]= 1426685652;
assign addr[22648]= 1368621831;
assign addr[22649]= 1308821808;
assign addr[22650]= 1247361445;
assign addr[22651]= 1184318708;
assign addr[22652]= 1119773573;
assign addr[22653]= 1053807919;
assign addr[22654]= 986505429;
assign addr[22655]= 917951481;
assign addr[22656]= 848233042;
assign addr[22657]= 777438554;
assign addr[22658]= 705657826;
assign addr[22659]= 632981917;
assign addr[22660]= 559503022;
assign addr[22661]= 485314355;
assign addr[22662]= 410510029;
assign addr[22663]= 335184940;
assign addr[22664]= 259434643;
assign addr[22665]= 183355234;
assign addr[22666]= 107043224;
assign addr[22667]= 30595422;
assign addr[22668]= -45891193;
assign addr[22669]= -122319591;
assign addr[22670]= -198592817;
assign addr[22671]= -274614114;
assign addr[22672]= -350287041;
assign addr[22673]= -425515602;
assign addr[22674]= -500204365;
assign addr[22675]= -574258580;
assign addr[22676]= -647584304;
assign addr[22677]= -720088517;
assign addr[22678]= -791679244;
assign addr[22679]= -862265664;
assign addr[22680]= -931758235;
assign addr[22681]= -1000068799;
assign addr[22682]= -1067110699;
assign addr[22683]= -1132798888;
assign addr[22684]= -1197050035;
assign addr[22685]= -1259782632;
assign addr[22686]= -1320917099;
assign addr[22687]= -1380375881;
assign addr[22688]= -1438083551;
assign addr[22689]= -1493966902;
assign addr[22690]= -1547955041;
assign addr[22691]= -1599979481;
assign addr[22692]= -1649974225;
assign addr[22693]= -1697875851;
assign addr[22694]= -1743623590;
assign addr[22695]= -1787159411;
assign addr[22696]= -1828428082;
assign addr[22697]= -1867377253;
assign addr[22698]= -1903957513;
assign addr[22699]= -1938122457;
assign addr[22700]= -1969828744;
assign addr[22701]= -1999036154;
assign addr[22702]= -2025707632;
assign addr[22703]= -2049809346;
assign addr[22704]= -2071310720;
assign addr[22705]= -2090184478;
assign addr[22706]= -2106406677;
assign addr[22707]= -2119956737;
assign addr[22708]= -2130817471;
assign addr[22709]= -2138975100;
assign addr[22710]= -2144419275;
assign addr[22711]= -2147143090;
assign addr[22712]= -2147143090;
assign addr[22713]= -2144419275;
assign addr[22714]= -2138975100;
assign addr[22715]= -2130817471;
assign addr[22716]= -2119956737;
assign addr[22717]= -2106406677;
assign addr[22718]= -2090184478;
assign addr[22719]= -2071310720;
assign addr[22720]= -2049809346;
assign addr[22721]= -2025707632;
assign addr[22722]= -1999036154;
assign addr[22723]= -1969828744;
assign addr[22724]= -1938122457;
assign addr[22725]= -1903957513;
assign addr[22726]= -1867377253;
assign addr[22727]= -1828428082;
assign addr[22728]= -1787159411;
assign addr[22729]= -1743623590;
assign addr[22730]= -1697875851;
assign addr[22731]= -1649974225;
assign addr[22732]= -1599979481;
assign addr[22733]= -1547955041;
assign addr[22734]= -1493966902;
assign addr[22735]= -1438083551;
assign addr[22736]= -1380375881;
assign addr[22737]= -1320917099;
assign addr[22738]= -1259782632;
assign addr[22739]= -1197050035;
assign addr[22740]= -1132798888;
assign addr[22741]= -1067110699;
assign addr[22742]= -1000068799;
assign addr[22743]= -931758235;
assign addr[22744]= -862265664;
assign addr[22745]= -791679244;
assign addr[22746]= -720088517;
assign addr[22747]= -647584304;
assign addr[22748]= -574258580;
assign addr[22749]= -500204365;
assign addr[22750]= -425515602;
assign addr[22751]= -350287041;
assign addr[22752]= -274614114;
assign addr[22753]= -198592817;
assign addr[22754]= -122319591;
assign addr[22755]= -45891193;
assign addr[22756]= 30595422;
assign addr[22757]= 107043224;
assign addr[22758]= 183355234;
assign addr[22759]= 259434643;
assign addr[22760]= 335184940;
assign addr[22761]= 410510029;
assign addr[22762]= 485314355;
assign addr[22763]= 559503022;
assign addr[22764]= 632981917;
assign addr[22765]= 705657826;
assign addr[22766]= 777438554;
assign addr[22767]= 848233042;
assign addr[22768]= 917951481;
assign addr[22769]= 986505429;
assign addr[22770]= 1053807919;
assign addr[22771]= 1119773573;
assign addr[22772]= 1184318708;
assign addr[22773]= 1247361445;
assign addr[22774]= 1308821808;
assign addr[22775]= 1368621831;
assign addr[22776]= 1426685652;
assign addr[22777]= 1482939614;
assign addr[22778]= 1537312353;
assign addr[22779]= 1589734894;
assign addr[22780]= 1640140734;
assign addr[22781]= 1688465931;
assign addr[22782]= 1734649179;
assign addr[22783]= 1778631892;
assign addr[22784]= 1820358275;
assign addr[22785]= 1859775393;
assign addr[22786]= 1896833245;
assign addr[22787]= 1931484818;
assign addr[22788]= 1963686155;
assign addr[22789]= 1993396407;
assign addr[22790]= 2020577882;
assign addr[22791]= 2045196100;
assign addr[22792]= 2067219829;
assign addr[22793]= 2086621133;
assign addr[22794]= 2103375398;
assign addr[22795]= 2117461370;
assign addr[22796]= 2128861181;
assign addr[22797]= 2137560369;
assign addr[22798]= 2143547897;
assign addr[22799]= 2146816171;
assign addr[22800]= 2147361045;
assign addr[22801]= 2145181827;
assign addr[22802]= 2140281282;
assign addr[22803]= 2132665626;
assign addr[22804]= 2122344521;
assign addr[22805]= 2109331059;
assign addr[22806]= 2093641749;
assign addr[22807]= 2075296495;
assign addr[22808]= 2054318569;
assign addr[22809]= 2030734582;
assign addr[22810]= 2004574453;
assign addr[22811]= 1975871368;
assign addr[22812]= 1944661739;
assign addr[22813]= 1910985158;
assign addr[22814]= 1874884346;
assign addr[22815]= 1836405100;
assign addr[22816]= 1795596234;
assign addr[22817]= 1752509516;
assign addr[22818]= 1707199606;
assign addr[22819]= 1659723983;
assign addr[22820]= 1610142873;
assign addr[22821]= 1558519173;
assign addr[22822]= 1504918373;
assign addr[22823]= 1449408469;
assign addr[22824]= 1392059879;
assign addr[22825]= 1332945355;
assign addr[22826]= 1272139887;
assign addr[22827]= 1209720613;
assign addr[22828]= 1145766716;
assign addr[22829]= 1080359326;
assign addr[22830]= 1013581418;
assign addr[22831]= 945517704;
assign addr[22832]= 876254528;
assign addr[22833]= 805879757;
assign addr[22834]= 734482665;
assign addr[22835]= 662153826;
assign addr[22836]= 588984994;
assign addr[22837]= 515068990;
assign addr[22838]= 440499581;
assign addr[22839]= 365371365;
assign addr[22840]= 289779648;
assign addr[22841]= 213820322;
assign addr[22842]= 137589750;
assign addr[22843]= 61184634;
assign addr[22844]= -15298099;
assign addr[22845]= -91761426;
assign addr[22846]= -168108346;
assign addr[22847]= -244242007;
assign addr[22848]= -320065829;
assign addr[22849]= -395483624;
assign addr[22850]= -470399716;
assign addr[22851]= -544719071;
assign addr[22852]= -618347408;
assign addr[22853]= -691191324;
assign addr[22854]= -763158411;
assign addr[22855]= -834157373;
assign addr[22856]= -904098143;
assign addr[22857]= -972891995;
assign addr[22858]= -1040451659;
assign addr[22859]= -1106691431;
assign addr[22860]= -1171527280;
assign addr[22861]= -1234876957;
assign addr[22862]= -1296660098;
assign addr[22863]= -1356798326;
assign addr[22864]= -1415215352;
assign addr[22865]= -1471837070;
assign addr[22866]= -1526591649;
assign addr[22867]= -1579409630;
assign addr[22868]= -1630224009;
assign addr[22869]= -1678970324;
assign addr[22870]= -1725586737;
assign addr[22871]= -1770014111;
assign addr[22872]= -1812196087;
assign addr[22873]= -1852079154;
assign addr[22874]= -1889612716;
assign addr[22875]= -1924749160;
assign addr[22876]= -1957443913;
assign addr[22877]= -1987655498;
assign addr[22878]= -2015345591;
assign addr[22879]= -2040479063;
assign addr[22880]= -2063024031;
assign addr[22881]= -2082951896;
assign addr[22882]= -2100237377;
assign addr[22883]= -2114858546;
assign addr[22884]= -2126796855;
assign addr[22885]= -2136037160;
assign addr[22886]= -2142567738;
assign addr[22887]= -2146380306;
assign addr[22888]= -2147470025;
assign addr[22889]= -2145835515;
assign addr[22890]= -2141478848;
assign addr[22891]= -2134405552;
assign addr[22892]= -2124624598;
assign addr[22893]= -2112148396;
assign addr[22894]= -2096992772;
assign addr[22895]= -2079176953;
assign addr[22896]= -2058723538;
assign addr[22897]= -2035658475;
assign addr[22898]= -2010011024;
assign addr[22899]= -1981813720;
assign addr[22900]= -1951102334;
assign addr[22901]= -1917915825;
assign addr[22902]= -1882296293;
assign addr[22903]= -1844288924;
assign addr[22904]= -1803941934;
assign addr[22905]= -1761306505;
assign addr[22906]= -1716436725;
assign addr[22907]= -1669389513;
assign addr[22908]= -1620224553;
assign addr[22909]= -1569004214;
assign addr[22910]= -1515793473;
assign addr[22911]= -1460659832;
assign addr[22912]= -1403673233;
assign addr[22913]= -1344905966;
assign addr[22914]= -1284432584;
assign addr[22915]= -1222329801;
assign addr[22916]= -1158676398;
assign addr[22917]= -1093553126;
assign addr[22918]= -1027042599;
assign addr[22919]= -959229189;
assign addr[22920]= -890198924;
assign addr[22921]= -820039373;
assign addr[22922]= -748839539;
assign addr[22923]= -676689746;
assign addr[22924]= -603681519;
assign addr[22925]= -529907477;
assign addr[22926]= -455461206;
assign addr[22927]= -380437148;
assign addr[22928]= -304930476;
assign addr[22929]= -229036977;
assign addr[22930]= -152852926;
assign addr[22931]= -76474970;
assign addr[22932]= 0;
assign addr[22933]= 76474970;
assign addr[22934]= 152852926;
assign addr[22935]= 229036977;
assign addr[22936]= 304930476;
assign addr[22937]= 380437148;
assign addr[22938]= 455461206;
assign addr[22939]= 529907477;
assign addr[22940]= 603681519;
assign addr[22941]= 676689746;
assign addr[22942]= 748839539;
assign addr[22943]= 820039373;
assign addr[22944]= 890198924;
assign addr[22945]= 959229189;
assign addr[22946]= 1027042599;
assign addr[22947]= 1093553126;
assign addr[22948]= 1158676398;
assign addr[22949]= 1222329801;
assign addr[22950]= 1284432584;
assign addr[22951]= 1344905966;
assign addr[22952]= 1403673233;
assign addr[22953]= 1460659832;
assign addr[22954]= 1515793473;
assign addr[22955]= 1569004214;
assign addr[22956]= 1620224553;
assign addr[22957]= 1669389513;
assign addr[22958]= 1716436725;
assign addr[22959]= 1761306505;
assign addr[22960]= 1803941934;
assign addr[22961]= 1844288924;
assign addr[22962]= 1882296293;
assign addr[22963]= 1917915825;
assign addr[22964]= 1951102334;
assign addr[22965]= 1981813720;
assign addr[22966]= 2010011024;
assign addr[22967]= 2035658475;
assign addr[22968]= 2058723538;
assign addr[22969]= 2079176953;
assign addr[22970]= 2096992772;
assign addr[22971]= 2112148396;
assign addr[22972]= 2124624598;
assign addr[22973]= 2134405552;
assign addr[22974]= 2141478848;
assign addr[22975]= 2145835515;
assign addr[22976]= 2147470025;
assign addr[22977]= 2146380306;
assign addr[22978]= 2142567738;
assign addr[22979]= 2136037160;
assign addr[22980]= 2126796855;
assign addr[22981]= 2114858546;
assign addr[22982]= 2100237377;
assign addr[22983]= 2082951896;
assign addr[22984]= 2063024031;
assign addr[22985]= 2040479063;
assign addr[22986]= 2015345591;
assign addr[22987]= 1987655498;
assign addr[22988]= 1957443913;
assign addr[22989]= 1924749160;
assign addr[22990]= 1889612716;
assign addr[22991]= 1852079154;
assign addr[22992]= 1812196087;
assign addr[22993]= 1770014111;
assign addr[22994]= 1725586737;
assign addr[22995]= 1678970324;
assign addr[22996]= 1630224009;
assign addr[22997]= 1579409630;
assign addr[22998]= 1526591649;
assign addr[22999]= 1471837070;
assign addr[23000]= 1415215352;
assign addr[23001]= 1356798326;
assign addr[23002]= 1296660098;
assign addr[23003]= 1234876957;
assign addr[23004]= 1171527280;
assign addr[23005]= 1106691431;
assign addr[23006]= 1040451659;
assign addr[23007]= 972891995;
assign addr[23008]= 904098143;
assign addr[23009]= 834157373;
assign addr[23010]= 763158411;
assign addr[23011]= 691191324;
assign addr[23012]= 618347408;
assign addr[23013]= 544719071;
assign addr[23014]= 470399716;
assign addr[23015]= 395483624;
assign addr[23016]= 320065829;
assign addr[23017]= 244242007;
assign addr[23018]= 168108346;
assign addr[23019]= 91761426;
assign addr[23020]= 15298099;
assign addr[23021]= -61184634;
assign addr[23022]= -137589750;
assign addr[23023]= -213820322;
assign addr[23024]= -289779648;
assign addr[23025]= -365371365;
assign addr[23026]= -440499581;
assign addr[23027]= -515068990;
assign addr[23028]= -588984994;
assign addr[23029]= -662153826;
assign addr[23030]= -734482665;
assign addr[23031]= -805879757;
assign addr[23032]= -876254528;
assign addr[23033]= -945517704;
assign addr[23034]= -1013581418;
assign addr[23035]= -1080359326;
assign addr[23036]= -1145766716;
assign addr[23037]= -1209720613;
assign addr[23038]= -1272139887;
assign addr[23039]= -1332945355;
assign addr[23040]= -1392059879;
assign addr[23041]= -1449408469;
assign addr[23042]= -1504918373;
assign addr[23043]= -1558519173;
assign addr[23044]= -1610142873;
assign addr[23045]= -1659723983;
assign addr[23046]= -1707199606;
assign addr[23047]= -1752509516;
assign addr[23048]= -1795596234;
assign addr[23049]= -1836405100;
assign addr[23050]= -1874884346;
assign addr[23051]= -1910985158;
assign addr[23052]= -1944661739;
assign addr[23053]= -1975871368;
assign addr[23054]= -2004574453;
assign addr[23055]= -2030734582;
assign addr[23056]= -2054318569;
assign addr[23057]= -2075296495;
assign addr[23058]= -2093641749;
assign addr[23059]= -2109331059;
assign addr[23060]= -2122344521;
assign addr[23061]= -2132665626;
assign addr[23062]= -2140281282;
assign addr[23063]= -2145181827;
assign addr[23064]= -2147361045;
assign addr[23065]= -2146816171;
assign addr[23066]= -2143547897;
assign addr[23067]= -2137560369;
assign addr[23068]= -2128861181;
assign addr[23069]= -2117461370;
assign addr[23070]= -2103375398;
assign addr[23071]= -2086621133;
assign addr[23072]= -2067219829;
assign addr[23073]= -2045196100;
assign addr[23074]= -2020577882;
assign addr[23075]= -1993396407;
assign addr[23076]= -1963686155;
assign addr[23077]= -1931484818;
assign addr[23078]= -1896833245;
assign addr[23079]= -1859775393;
assign addr[23080]= -1820358275;
assign addr[23081]= -1778631892;
assign addr[23082]= -1734649179;
assign addr[23083]= -1688465931;
assign addr[23084]= -1640140734;
assign addr[23085]= -1589734894;
assign addr[23086]= -1537312353;
assign addr[23087]= -1482939614;
assign addr[23088]= -1426685652;
assign addr[23089]= -1368621831;
assign addr[23090]= -1308821808;
assign addr[23091]= -1247361445;
assign addr[23092]= -1184318708;
assign addr[23093]= -1119773573;
assign addr[23094]= -1053807919;
assign addr[23095]= -986505429;
assign addr[23096]= -917951481;
assign addr[23097]= -848233042;
assign addr[23098]= -777438554;
assign addr[23099]= -705657826;
assign addr[23100]= -632981917;
assign addr[23101]= -559503022;
assign addr[23102]= -485314355;
assign addr[23103]= -410510029;
assign addr[23104]= -335184940;
assign addr[23105]= -259434643;
assign addr[23106]= -183355234;
assign addr[23107]= -107043224;
assign addr[23108]= -30595422;
assign addr[23109]= 45891193;
assign addr[23110]= 122319591;
assign addr[23111]= 198592817;
assign addr[23112]= 274614114;
assign addr[23113]= 350287041;
assign addr[23114]= 425515602;
assign addr[23115]= 500204365;
assign addr[23116]= 574258580;
assign addr[23117]= 647584304;
assign addr[23118]= 720088517;
assign addr[23119]= 791679244;
assign addr[23120]= 862265664;
assign addr[23121]= 931758235;
assign addr[23122]= 1000068799;
assign addr[23123]= 1067110699;
assign addr[23124]= 1132798888;
assign addr[23125]= 1197050035;
assign addr[23126]= 1259782632;
assign addr[23127]= 1320917099;
assign addr[23128]= 1380375881;
assign addr[23129]= 1438083551;
assign addr[23130]= 1493966902;
assign addr[23131]= 1547955041;
assign addr[23132]= 1599979481;
assign addr[23133]= 1649974225;
assign addr[23134]= 1697875851;
assign addr[23135]= 1743623590;
assign addr[23136]= 1787159411;
assign addr[23137]= 1828428082;
assign addr[23138]= 1867377253;
assign addr[23139]= 1903957513;
assign addr[23140]= 1938122457;
assign addr[23141]= 1969828744;
assign addr[23142]= 1999036154;
assign addr[23143]= 2025707632;
assign addr[23144]= 2049809346;
assign addr[23145]= 2071310720;
assign addr[23146]= 2090184478;
assign addr[23147]= 2106406677;
assign addr[23148]= 2119956737;
assign addr[23149]= 2130817471;
assign addr[23150]= 2138975100;
assign addr[23151]= 2144419275;
assign addr[23152]= 2147143090;
assign addr[23153]= 2147143090;
assign addr[23154]= 2144419275;
assign addr[23155]= 2138975100;
assign addr[23156]= 2130817471;
assign addr[23157]= 2119956737;
assign addr[23158]= 2106406677;
assign addr[23159]= 2090184478;
assign addr[23160]= 2071310720;
assign addr[23161]= 2049809346;
assign addr[23162]= 2025707632;
assign addr[23163]= 1999036154;
assign addr[23164]= 1969828744;
assign addr[23165]= 1938122457;
assign addr[23166]= 1903957513;
assign addr[23167]= 1867377253;
assign addr[23168]= 1828428082;
assign addr[23169]= 1787159411;
assign addr[23170]= 1743623590;
assign addr[23171]= 1697875851;
assign addr[23172]= 1649974225;
assign addr[23173]= 1599979481;
assign addr[23174]= 1547955041;
assign addr[23175]= 1493966902;
assign addr[23176]= 1438083551;
assign addr[23177]= 1380375881;
assign addr[23178]= 1320917099;
assign addr[23179]= 1259782632;
assign addr[23180]= 1197050035;
assign addr[23181]= 1132798888;
assign addr[23182]= 1067110699;
assign addr[23183]= 1000068799;
assign addr[23184]= 931758235;
assign addr[23185]= 862265664;
assign addr[23186]= 791679244;
assign addr[23187]= 720088517;
assign addr[23188]= 647584304;
assign addr[23189]= 574258580;
assign addr[23190]= 500204365;
assign addr[23191]= 425515602;
assign addr[23192]= 350287041;
assign addr[23193]= 274614114;
assign addr[23194]= 198592817;
assign addr[23195]= 122319591;
assign addr[23196]= 45891193;
assign addr[23197]= -30595422;
assign addr[23198]= -107043224;
assign addr[23199]= -183355234;
assign addr[23200]= -259434643;
assign addr[23201]= -335184940;
assign addr[23202]= -410510029;
assign addr[23203]= -485314355;
assign addr[23204]= -559503022;
assign addr[23205]= -632981917;
assign addr[23206]= -705657826;
assign addr[23207]= -777438554;
assign addr[23208]= -848233042;
assign addr[23209]= -917951481;
assign addr[23210]= -986505429;
assign addr[23211]= -1053807919;
assign addr[23212]= -1119773573;
assign addr[23213]= -1184318708;
assign addr[23214]= -1247361445;
assign addr[23215]= -1308821808;
assign addr[23216]= -1368621831;
assign addr[23217]= -1426685652;
assign addr[23218]= -1482939614;
assign addr[23219]= -1537312353;
assign addr[23220]= -1589734894;
assign addr[23221]= -1640140734;
assign addr[23222]= -1688465931;
assign addr[23223]= -1734649179;
assign addr[23224]= -1778631892;
assign addr[23225]= -1820358275;
assign addr[23226]= -1859775393;
assign addr[23227]= -1896833245;
assign addr[23228]= -1931484818;
assign addr[23229]= -1963686155;
assign addr[23230]= -1993396407;
assign addr[23231]= -2020577882;
assign addr[23232]= -2045196100;
assign addr[23233]= -2067219829;
assign addr[23234]= -2086621133;
assign addr[23235]= -2103375398;
assign addr[23236]= -2117461370;
assign addr[23237]= -2128861181;
assign addr[23238]= -2137560369;
assign addr[23239]= -2143547897;
assign addr[23240]= -2146816171;
assign addr[23241]= -2147361045;
assign addr[23242]= -2145181827;
assign addr[23243]= -2140281282;
assign addr[23244]= -2132665626;
assign addr[23245]= -2122344521;
assign addr[23246]= -2109331059;
assign addr[23247]= -2093641749;
assign addr[23248]= -2075296495;
assign addr[23249]= -2054318569;
assign addr[23250]= -2030734582;
assign addr[23251]= -2004574453;
assign addr[23252]= -1975871368;
assign addr[23253]= -1944661739;
assign addr[23254]= -1910985158;
assign addr[23255]= -1874884346;
assign addr[23256]= -1836405100;
assign addr[23257]= -1795596234;
assign addr[23258]= -1752509516;
assign addr[23259]= -1707199606;
assign addr[23260]= -1659723983;
assign addr[23261]= -1610142873;
assign addr[23262]= -1558519173;
assign addr[23263]= -1504918373;
assign addr[23264]= -1449408469;
assign addr[23265]= -1392059879;
assign addr[23266]= -1332945355;
assign addr[23267]= -1272139887;
assign addr[23268]= -1209720613;
assign addr[23269]= -1145766716;
assign addr[23270]= -1080359326;
assign addr[23271]= -1013581418;
assign addr[23272]= -945517704;
assign addr[23273]= -876254528;
assign addr[23274]= -805879757;
assign addr[23275]= -734482665;
assign addr[23276]= -662153826;
assign addr[23277]= -588984994;
assign addr[23278]= -515068990;
assign addr[23279]= -440499581;
assign addr[23280]= -365371365;
assign addr[23281]= -289779648;
assign addr[23282]= -213820322;
assign addr[23283]= -137589750;
assign addr[23284]= -61184634;
assign addr[23285]= 15298099;
assign addr[23286]= 91761426;
assign addr[23287]= 168108346;
assign addr[23288]= 244242007;
assign addr[23289]= 320065829;
assign addr[23290]= 395483624;
assign addr[23291]= 470399716;
assign addr[23292]= 544719071;
assign addr[23293]= 618347408;
assign addr[23294]= 691191324;
assign addr[23295]= 763158411;
assign addr[23296]= 834157373;
assign addr[23297]= 904098143;
assign addr[23298]= 972891995;
assign addr[23299]= 1040451659;
assign addr[23300]= 1106691431;
assign addr[23301]= 1171527280;
assign addr[23302]= 1234876957;
assign addr[23303]= 1296660098;
assign addr[23304]= 1356798326;
assign addr[23305]= 1415215352;
assign addr[23306]= 1471837070;
assign addr[23307]= 1526591649;
assign addr[23308]= 1579409630;
assign addr[23309]= 1630224009;
assign addr[23310]= 1678970324;
assign addr[23311]= 1725586737;
assign addr[23312]= 1770014111;
assign addr[23313]= 1812196087;
assign addr[23314]= 1852079154;
assign addr[23315]= 1889612716;
assign addr[23316]= 1924749160;
assign addr[23317]= 1957443913;
assign addr[23318]= 1987655498;
assign addr[23319]= 2015345591;
assign addr[23320]= 2040479063;
assign addr[23321]= 2063024031;
assign addr[23322]= 2082951896;
assign addr[23323]= 2100237377;
assign addr[23324]= 2114858546;
assign addr[23325]= 2126796855;
assign addr[23326]= 2136037160;
assign addr[23327]= 2142567738;
assign addr[23328]= 2146380306;
assign addr[23329]= 2147470025;
assign addr[23330]= 2145835515;
assign addr[23331]= 2141478848;
assign addr[23332]= 2134405552;
assign addr[23333]= 2124624598;
assign addr[23334]= 2112148396;
assign addr[23335]= 2096992772;
assign addr[23336]= 2079176953;
assign addr[23337]= 2058723538;
assign addr[23338]= 2035658475;
assign addr[23339]= 2010011024;
assign addr[23340]= 1981813720;
assign addr[23341]= 1951102334;
assign addr[23342]= 1917915825;
assign addr[23343]= 1882296293;
assign addr[23344]= 1844288924;
assign addr[23345]= 1803941934;
assign addr[23346]= 1761306505;
assign addr[23347]= 1716436725;
assign addr[23348]= 1669389513;
assign addr[23349]= 1620224553;
assign addr[23350]= 1569004214;
assign addr[23351]= 1515793473;
assign addr[23352]= 1460659832;
assign addr[23353]= 1403673233;
assign addr[23354]= 1344905966;
assign addr[23355]= 1284432584;
assign addr[23356]= 1222329801;
assign addr[23357]= 1158676398;
assign addr[23358]= 1093553126;
assign addr[23359]= 1027042599;
assign addr[23360]= 959229189;
assign addr[23361]= 890198924;
assign addr[23362]= 820039373;
assign addr[23363]= 748839539;
assign addr[23364]= 676689746;
assign addr[23365]= 603681519;
assign addr[23366]= 529907477;
assign addr[23367]= 455461206;
assign addr[23368]= 380437148;
assign addr[23369]= 304930476;
assign addr[23370]= 229036977;
assign addr[23371]= 152852926;
assign addr[23372]= 76474970;
assign addr[23373]= 0;
assign addr[23374]= -76474970;
assign addr[23375]= -152852926;
assign addr[23376]= -229036977;
assign addr[23377]= -304930476;
assign addr[23378]= -380437148;
assign addr[23379]= -455461206;
assign addr[23380]= -529907477;
assign addr[23381]= -603681519;
assign addr[23382]= -676689746;
assign addr[23383]= -748839539;
assign addr[23384]= -820039373;
assign addr[23385]= -890198924;
assign addr[23386]= -959229189;
assign addr[23387]= -1027042599;
assign addr[23388]= -1093553126;
assign addr[23389]= -1158676398;
assign addr[23390]= -1222329801;
assign addr[23391]= -1284432584;
assign addr[23392]= -1344905966;
assign addr[23393]= -1403673233;
assign addr[23394]= -1460659832;
assign addr[23395]= -1515793473;
assign addr[23396]= -1569004214;
assign addr[23397]= -1620224553;
assign addr[23398]= -1669389513;
assign addr[23399]= -1716436725;
assign addr[23400]= -1761306505;
assign addr[23401]= -1803941934;
assign addr[23402]= -1844288924;
assign addr[23403]= -1882296293;
assign addr[23404]= -1917915825;
assign addr[23405]= -1951102334;
assign addr[23406]= -1981813720;
assign addr[23407]= -2010011024;
assign addr[23408]= -2035658475;
assign addr[23409]= -2058723538;
assign addr[23410]= -2079176953;
assign addr[23411]= -2096992772;
assign addr[23412]= -2112148396;
assign addr[23413]= -2124624598;
assign addr[23414]= -2134405552;
assign addr[23415]= -2141478848;
assign addr[23416]= -2145835515;
assign addr[23417]= -2147470025;
assign addr[23418]= -2146380306;
assign addr[23419]= -2142567738;
assign addr[23420]= -2136037160;
assign addr[23421]= -2126796855;
assign addr[23422]= -2114858546;
assign addr[23423]= -2100237377;
assign addr[23424]= -2082951896;
assign addr[23425]= -2063024031;
assign addr[23426]= -2040479063;
assign addr[23427]= -2015345591;
assign addr[23428]= -1987655498;
assign addr[23429]= -1957443913;
assign addr[23430]= -1924749160;
assign addr[23431]= -1889612716;
assign addr[23432]= -1852079154;
assign addr[23433]= -1812196087;
assign addr[23434]= -1770014111;
assign addr[23435]= -1725586737;
assign addr[23436]= -1678970324;
assign addr[23437]= -1630224009;
assign addr[23438]= -1579409630;
assign addr[23439]= -1526591649;
assign addr[23440]= -1471837070;
assign addr[23441]= -1415215352;
assign addr[23442]= -1356798326;
assign addr[23443]= -1296660098;
assign addr[23444]= -1234876957;
assign addr[23445]= -1171527280;
assign addr[23446]= -1106691431;
assign addr[23447]= -1040451659;
assign addr[23448]= -972891995;
assign addr[23449]= -904098143;
assign addr[23450]= -834157373;
assign addr[23451]= -763158411;
assign addr[23452]= -691191324;
assign addr[23453]= -618347408;
assign addr[23454]= -544719071;
assign addr[23455]= -470399716;
assign addr[23456]= -395483624;
assign addr[23457]= -320065829;
assign addr[23458]= -244242007;
assign addr[23459]= -168108346;
assign addr[23460]= -91761426;
assign addr[23461]= -15298099;
assign addr[23462]= 61184634;
assign addr[23463]= 137589750;
assign addr[23464]= 213820322;
assign addr[23465]= 289779648;
assign addr[23466]= 365371365;
assign addr[23467]= 440499581;
assign addr[23468]= 515068990;
assign addr[23469]= 588984994;
assign addr[23470]= 662153826;
assign addr[23471]= 734482665;
assign addr[23472]= 805879757;
assign addr[23473]= 876254528;
assign addr[23474]= 945517704;
assign addr[23475]= 1013581418;
assign addr[23476]= 1080359326;
assign addr[23477]= 1145766716;
assign addr[23478]= 1209720613;
assign addr[23479]= 1272139887;
assign addr[23480]= 1332945355;
assign addr[23481]= 1392059879;
assign addr[23482]= 1449408469;
assign addr[23483]= 1504918373;
assign addr[23484]= 1558519173;
assign addr[23485]= 1610142873;
assign addr[23486]= 1659723983;
assign addr[23487]= 1707199606;
assign addr[23488]= 1752509516;
assign addr[23489]= 1795596234;
assign addr[23490]= 1836405100;
assign addr[23491]= 1874884346;
assign addr[23492]= 1910985158;
assign addr[23493]= 1944661739;
assign addr[23494]= 1975871368;
assign addr[23495]= 2004574453;
assign addr[23496]= 2030734582;
assign addr[23497]= 2054318569;
assign addr[23498]= 2075296495;
assign addr[23499]= 2093641749;
assign addr[23500]= 2109331059;
assign addr[23501]= 2122344521;
assign addr[23502]= 2132665626;
assign addr[23503]= 2140281282;
assign addr[23504]= 2145181827;
assign addr[23505]= 2147361045;
assign addr[23506]= 2146816171;
assign addr[23507]= 2143547897;
assign addr[23508]= 2137560369;
assign addr[23509]= 2128861181;
assign addr[23510]= 2117461370;
assign addr[23511]= 2103375398;
assign addr[23512]= 2086621133;
assign addr[23513]= 2067219829;
assign addr[23514]= 2045196100;
assign addr[23515]= 2020577882;
assign addr[23516]= 1993396407;
assign addr[23517]= 1963686155;
assign addr[23518]= 1931484818;
assign addr[23519]= 1896833245;
assign addr[23520]= 1859775393;
assign addr[23521]= 1820358275;
assign addr[23522]= 1778631892;
assign addr[23523]= 1734649179;
assign addr[23524]= 1688465931;
assign addr[23525]= 1640140734;
assign addr[23526]= 1589734894;
assign addr[23527]= 1537312353;
assign addr[23528]= 1482939614;
assign addr[23529]= 1426685652;
assign addr[23530]= 1368621831;
assign addr[23531]= 1308821808;
assign addr[23532]= 1247361445;
assign addr[23533]= 1184318708;
assign addr[23534]= 1119773573;
assign addr[23535]= 1053807919;
assign addr[23536]= 986505429;
assign addr[23537]= 917951481;
assign addr[23538]= 848233042;
assign addr[23539]= 777438554;
assign addr[23540]= 705657826;
assign addr[23541]= 632981917;
assign addr[23542]= 559503022;
assign addr[23543]= 485314355;
assign addr[23544]= 410510029;
assign addr[23545]= 335184940;
assign addr[23546]= 259434643;
assign addr[23547]= 183355234;
assign addr[23548]= 107043224;
assign addr[23549]= 30595422;
assign addr[23550]= -45891193;
assign addr[23551]= -122319591;
assign addr[23552]= -198592817;
assign addr[23553]= -274614114;
assign addr[23554]= -350287041;
assign addr[23555]= -425515602;
assign addr[23556]= -500204365;
assign addr[23557]= -574258580;
assign addr[23558]= -647584304;
assign addr[23559]= -720088517;
assign addr[23560]= -791679244;
assign addr[23561]= -862265664;
assign addr[23562]= -931758235;
assign addr[23563]= -1000068799;
assign addr[23564]= -1067110699;
assign addr[23565]= -1132798888;
assign addr[23566]= -1197050035;
assign addr[23567]= -1259782632;
assign addr[23568]= -1320917099;
assign addr[23569]= -1380375881;
assign addr[23570]= -1438083551;
assign addr[23571]= -1493966902;
assign addr[23572]= -1547955041;
assign addr[23573]= -1599979481;
assign addr[23574]= -1649974225;
assign addr[23575]= -1697875851;
assign addr[23576]= -1743623590;
assign addr[23577]= -1787159411;
assign addr[23578]= -1828428082;
assign addr[23579]= -1867377253;
assign addr[23580]= -1903957513;
assign addr[23581]= -1938122457;
assign addr[23582]= -1969828744;
assign addr[23583]= -1999036154;
assign addr[23584]= -2025707632;
assign addr[23585]= -2049809346;
assign addr[23586]= -2071310720;
assign addr[23587]= -2090184478;
assign addr[23588]= -2106406677;
assign addr[23589]= -2119956737;
assign addr[23590]= -2130817471;
assign addr[23591]= -2138975100;
assign addr[23592]= -2144419275;
assign addr[23593]= -2147143090;
assign addr[23594]= -2147143090;
assign addr[23595]= -2144419275;
assign addr[23596]= -2138975100;
assign addr[23597]= -2130817471;
assign addr[23598]= -2119956737;
assign addr[23599]= -2106406677;
assign addr[23600]= -2090184478;
assign addr[23601]= -2071310720;
assign addr[23602]= -2049809346;
assign addr[23603]= -2025707632;
assign addr[23604]= -1999036154;
assign addr[23605]= -1969828744;
assign addr[23606]= -1938122457;
assign addr[23607]= -1903957513;
assign addr[23608]= -1867377253;
assign addr[23609]= -1828428082;
assign addr[23610]= -1787159411;
assign addr[23611]= -1743623590;
assign addr[23612]= -1697875851;
assign addr[23613]= -1649974225;
assign addr[23614]= -1599979481;
assign addr[23615]= -1547955041;
assign addr[23616]= -1493966902;
assign addr[23617]= -1438083551;
assign addr[23618]= -1380375881;
assign addr[23619]= -1320917099;
assign addr[23620]= -1259782632;
assign addr[23621]= -1197050035;
assign addr[23622]= -1132798888;
assign addr[23623]= -1067110699;
assign addr[23624]= -1000068799;
assign addr[23625]= -931758235;
assign addr[23626]= -862265664;
assign addr[23627]= -791679244;
assign addr[23628]= -720088517;
assign addr[23629]= -647584304;
assign addr[23630]= -574258580;
assign addr[23631]= -500204365;
assign addr[23632]= -425515602;
assign addr[23633]= -350287041;
assign addr[23634]= -274614114;
assign addr[23635]= -198592817;
assign addr[23636]= -122319591;
assign addr[23637]= -45891193;
assign addr[23638]= 30595422;
assign addr[23639]= 107043224;
assign addr[23640]= 183355234;
assign addr[23641]= 259434643;
assign addr[23642]= 335184940;
assign addr[23643]= 410510029;
assign addr[23644]= 485314355;
assign addr[23645]= 559503022;
assign addr[23646]= 632981917;
assign addr[23647]= 705657826;
assign addr[23648]= 777438554;
assign addr[23649]= 848233042;
assign addr[23650]= 917951481;
assign addr[23651]= 986505429;
assign addr[23652]= 1053807919;
assign addr[23653]= 1119773573;
assign addr[23654]= 1184318708;
assign addr[23655]= 1247361445;
assign addr[23656]= 1308821808;
assign addr[23657]= 1368621831;
assign addr[23658]= 1426685652;
assign addr[23659]= 1482939614;
assign addr[23660]= 1537312353;
assign addr[23661]= 1589734894;
assign addr[23662]= 1640140734;
assign addr[23663]= 1688465931;
assign addr[23664]= 1734649179;
assign addr[23665]= 1778631892;
assign addr[23666]= 1820358275;
assign addr[23667]= 1859775393;
assign addr[23668]= 1896833245;
assign addr[23669]= 1931484818;
assign addr[23670]= 1963686155;
assign addr[23671]= 1993396407;
assign addr[23672]= 2020577882;
assign addr[23673]= 2045196100;
assign addr[23674]= 2067219829;
assign addr[23675]= 2086621133;
assign addr[23676]= 2103375398;
assign addr[23677]= 2117461370;
assign addr[23678]= 2128861181;
assign addr[23679]= 2137560369;
assign addr[23680]= 2143547897;
assign addr[23681]= 2146816171;
assign addr[23682]= 2147361045;
assign addr[23683]= 2145181827;
assign addr[23684]= 2140281282;
assign addr[23685]= 2132665626;
assign addr[23686]= 2122344521;
assign addr[23687]= 2109331059;
assign addr[23688]= 2093641749;
assign addr[23689]= 2075296495;
assign addr[23690]= 2054318569;
assign addr[23691]= 2030734582;
assign addr[23692]= 2004574453;
assign addr[23693]= 1975871368;
assign addr[23694]= 1944661739;
assign addr[23695]= 1910985158;
assign addr[23696]= 1874884346;
assign addr[23697]= 1836405100;
assign addr[23698]= 1795596234;
assign addr[23699]= 1752509516;
assign addr[23700]= 1707199606;
assign addr[23701]= 1659723983;
assign addr[23702]= 1610142873;
assign addr[23703]= 1558519173;
assign addr[23704]= 1504918373;
assign addr[23705]= 1449408469;
assign addr[23706]= 1392059879;
assign addr[23707]= 1332945355;
assign addr[23708]= 1272139887;
assign addr[23709]= 1209720613;
assign addr[23710]= 1145766716;
assign addr[23711]= 1080359326;
assign addr[23712]= 1013581418;
assign addr[23713]= 945517704;
assign addr[23714]= 876254528;
assign addr[23715]= 805879757;
assign addr[23716]= 734482665;
assign addr[23717]= 662153826;
assign addr[23718]= 588984994;
assign addr[23719]= 515068990;
assign addr[23720]= 440499581;
assign addr[23721]= 365371365;
assign addr[23722]= 289779648;
assign addr[23723]= 213820322;
assign addr[23724]= 137589750;
assign addr[23725]= 61184634;
assign addr[23726]= -15298099;
assign addr[23727]= -91761426;
assign addr[23728]= -168108346;
assign addr[23729]= -244242007;
assign addr[23730]= -320065829;
assign addr[23731]= -395483624;
assign addr[23732]= -470399716;
assign addr[23733]= -544719071;
assign addr[23734]= -618347408;
assign addr[23735]= -691191324;
assign addr[23736]= -763158411;
assign addr[23737]= -834157373;
assign addr[23738]= -904098143;
assign addr[23739]= -972891995;
assign addr[23740]= -1040451659;
assign addr[23741]= -1106691431;
assign addr[23742]= -1171527280;
assign addr[23743]= -1234876957;
assign addr[23744]= -1296660098;
assign addr[23745]= -1356798326;
assign addr[23746]= -1415215352;
assign addr[23747]= -1471837070;
assign addr[23748]= -1526591649;
assign addr[23749]= -1579409630;
assign addr[23750]= -1630224009;
assign addr[23751]= -1678970324;
assign addr[23752]= -1725586737;
assign addr[23753]= -1770014111;
assign addr[23754]= -1812196087;
assign addr[23755]= -1852079154;
assign addr[23756]= -1889612716;
assign addr[23757]= -1924749160;
assign addr[23758]= -1957443913;
assign addr[23759]= -1987655498;
assign addr[23760]= -2015345591;
assign addr[23761]= -2040479063;
assign addr[23762]= -2063024031;
assign addr[23763]= -2082951896;
assign addr[23764]= -2100237377;
assign addr[23765]= -2114858546;
assign addr[23766]= -2126796855;
assign addr[23767]= -2136037160;
assign addr[23768]= -2142567738;
assign addr[23769]= -2146380306;
assign addr[23770]= -2147470025;
assign addr[23771]= -2145835515;
assign addr[23772]= -2141478848;
assign addr[23773]= -2134405552;
assign addr[23774]= -2124624598;
assign addr[23775]= -2112148396;
assign addr[23776]= -2096992772;
assign addr[23777]= -2079176953;
assign addr[23778]= -2058723538;
assign addr[23779]= -2035658475;
assign addr[23780]= -2010011024;
assign addr[23781]= -1981813720;
assign addr[23782]= -1951102334;
assign addr[23783]= -1917915825;
assign addr[23784]= -1882296293;
assign addr[23785]= -1844288924;
assign addr[23786]= -1803941934;
assign addr[23787]= -1761306505;
assign addr[23788]= -1716436725;
assign addr[23789]= -1669389513;
assign addr[23790]= -1620224553;
assign addr[23791]= -1569004214;
assign addr[23792]= -1515793473;
assign addr[23793]= -1460659832;
assign addr[23794]= -1403673233;
assign addr[23795]= -1344905966;
assign addr[23796]= -1284432584;
assign addr[23797]= -1222329801;
assign addr[23798]= -1158676398;
assign addr[23799]= -1093553126;
assign addr[23800]= -1027042599;
assign addr[23801]= -959229189;
assign addr[23802]= -890198924;
assign addr[23803]= -820039373;
assign addr[23804]= -748839539;
assign addr[23805]= -676689746;
assign addr[23806]= -603681519;
assign addr[23807]= -529907477;
assign addr[23808]= -455461206;
assign addr[23809]= -380437148;
assign addr[23810]= -304930476;
assign addr[23811]= -229036977;
assign addr[23812]= -152852926;
assign addr[23813]= -76474970;
assign addr[23814]= 0;
assign addr[23815]= 76474970;
assign addr[23816]= 152852926;
assign addr[23817]= 229036977;
assign addr[23818]= 304930476;
assign addr[23819]= 380437148;
assign addr[23820]= 455461206;
assign addr[23821]= 529907477;
assign addr[23822]= 603681519;
assign addr[23823]= 676689746;
assign addr[23824]= 748839539;
assign addr[23825]= 820039373;
assign addr[23826]= 890198924;
assign addr[23827]= 959229189;
assign addr[23828]= 1027042599;
assign addr[23829]= 1093553126;
assign addr[23830]= 1158676398;
assign addr[23831]= 1222329801;
assign addr[23832]= 1284432584;
assign addr[23833]= 1344905966;
assign addr[23834]= 1403673233;
assign addr[23835]= 1460659832;
assign addr[23836]= 1515793473;
assign addr[23837]= 1569004214;
assign addr[23838]= 1620224553;
assign addr[23839]= 1669389513;
assign addr[23840]= 1716436725;
assign addr[23841]= 1761306505;
assign addr[23842]= 1803941934;
assign addr[23843]= 1844288924;
assign addr[23844]= 1882296293;
assign addr[23845]= 1917915825;
assign addr[23846]= 1951102334;
assign addr[23847]= 1981813720;
assign addr[23848]= 2010011024;
assign addr[23849]= 2035658475;
assign addr[23850]= 2058723538;
assign addr[23851]= 2079176953;
assign addr[23852]= 2096992772;
assign addr[23853]= 2112148396;
assign addr[23854]= 2124624598;
assign addr[23855]= 2134405552;
assign addr[23856]= 2141478848;
assign addr[23857]= 2145835515;
assign addr[23858]= 2147470025;
assign addr[23859]= 2146380306;
assign addr[23860]= 2142567738;
assign addr[23861]= 2136037160;
assign addr[23862]= 2126796855;
assign addr[23863]= 2114858546;
assign addr[23864]= 2100237377;
assign addr[23865]= 2082951896;
assign addr[23866]= 2063024031;
assign addr[23867]= 2040479063;
assign addr[23868]= 2015345591;
assign addr[23869]= 1987655498;
assign addr[23870]= 1957443913;
assign addr[23871]= 1924749160;
assign addr[23872]= 1889612716;
assign addr[23873]= 1852079154;
assign addr[23874]= 1812196087;
assign addr[23875]= 1770014111;
assign addr[23876]= 1725586737;
assign addr[23877]= 1678970324;
assign addr[23878]= 1630224009;
assign addr[23879]= 1579409630;
assign addr[23880]= 1526591649;
assign addr[23881]= 1471837070;
assign addr[23882]= 1415215352;
assign addr[23883]= 1356798326;
assign addr[23884]= 1296660098;
assign addr[23885]= 1234876957;
assign addr[23886]= 1171527280;
assign addr[23887]= 1106691431;
assign addr[23888]= 1040451659;
assign addr[23889]= 972891995;
assign addr[23890]= 904098143;
assign addr[23891]= 834157373;
assign addr[23892]= 763158411;
assign addr[23893]= 691191324;
assign addr[23894]= 618347408;
assign addr[23895]= 544719071;
assign addr[23896]= 470399716;
assign addr[23897]= 395483624;
assign addr[23898]= 320065829;
assign addr[23899]= 244242007;
assign addr[23900]= 168108346;
assign addr[23901]= 91761426;
assign addr[23902]= 15298099;
assign addr[23903]= -61184634;
assign addr[23904]= -137589750;
assign addr[23905]= -213820322;
assign addr[23906]= -289779648;
assign addr[23907]= -365371365;
assign addr[23908]= -440499581;
assign addr[23909]= -515068990;
assign addr[23910]= -588984994;
assign addr[23911]= -662153826;
assign addr[23912]= -734482665;
assign addr[23913]= -805879757;
assign addr[23914]= -876254528;
assign addr[23915]= -945517704;
assign addr[23916]= -1013581418;
assign addr[23917]= -1080359326;
assign addr[23918]= -1145766716;
assign addr[23919]= -1209720613;
assign addr[23920]= -1272139887;
assign addr[23921]= -1332945355;
assign addr[23922]= -1392059879;
assign addr[23923]= -1449408469;
assign addr[23924]= -1504918373;
assign addr[23925]= -1558519173;
assign addr[23926]= -1610142873;
assign addr[23927]= -1659723983;
assign addr[23928]= -1707199606;
assign addr[23929]= -1752509516;
assign addr[23930]= -1795596234;
assign addr[23931]= -1836405100;
assign addr[23932]= -1874884346;
assign addr[23933]= -1910985158;
assign addr[23934]= -1944661739;
assign addr[23935]= -1975871368;
assign addr[23936]= -2004574453;
assign addr[23937]= -2030734582;
assign addr[23938]= -2054318569;
assign addr[23939]= -2075296495;
assign addr[23940]= -2093641749;
assign addr[23941]= -2109331059;
assign addr[23942]= -2122344521;
assign addr[23943]= -2132665626;
assign addr[23944]= -2140281282;
assign addr[23945]= -2145181827;
assign addr[23946]= -2147361045;
assign addr[23947]= -2146816171;
assign addr[23948]= -2143547897;
assign addr[23949]= -2137560369;
assign addr[23950]= -2128861181;
assign addr[23951]= -2117461370;
assign addr[23952]= -2103375398;
assign addr[23953]= -2086621133;
assign addr[23954]= -2067219829;
assign addr[23955]= -2045196100;
assign addr[23956]= -2020577882;
assign addr[23957]= -1993396407;
assign addr[23958]= -1963686155;
assign addr[23959]= -1931484818;
assign addr[23960]= -1896833245;
assign addr[23961]= -1859775393;
assign addr[23962]= -1820358275;
assign addr[23963]= -1778631892;
assign addr[23964]= -1734649179;
assign addr[23965]= -1688465931;
assign addr[23966]= -1640140734;
assign addr[23967]= -1589734894;
assign addr[23968]= -1537312353;
assign addr[23969]= -1482939614;
assign addr[23970]= -1426685652;
assign addr[23971]= -1368621831;
assign addr[23972]= -1308821808;
assign addr[23973]= -1247361445;
assign addr[23974]= -1184318708;
assign addr[23975]= -1119773573;
assign addr[23976]= -1053807919;
assign addr[23977]= -986505429;
assign addr[23978]= -917951481;
assign addr[23979]= -848233042;
assign addr[23980]= -777438554;
assign addr[23981]= -705657826;
assign addr[23982]= -632981917;
assign addr[23983]= -559503022;
assign addr[23984]= -485314355;
assign addr[23985]= -410510029;
assign addr[23986]= -335184940;
assign addr[23987]= -259434643;
assign addr[23988]= -183355234;
assign addr[23989]= -107043224;
assign addr[23990]= -30595422;
assign addr[23991]= 45891193;
assign addr[23992]= 122319591;
assign addr[23993]= 198592817;
assign addr[23994]= 274614114;
assign addr[23995]= 350287041;
assign addr[23996]= 425515602;
assign addr[23997]= 500204365;
assign addr[23998]= 574258580;
assign addr[23999]= 647584304;
assign addr[24000]= 720088517;
assign addr[24001]= 791679244;
assign addr[24002]= 862265664;
assign addr[24003]= 931758235;
assign addr[24004]= 1000068799;
assign addr[24005]= 1067110699;
assign addr[24006]= 1132798888;
assign addr[24007]= 1197050035;
assign addr[24008]= 1259782632;
assign addr[24009]= 1320917099;
assign addr[24010]= 1380375881;
assign addr[24011]= 1438083551;
assign addr[24012]= 1493966902;
assign addr[24013]= 1547955041;
assign addr[24014]= 1599979481;
assign addr[24015]= 1649974225;
assign addr[24016]= 1697875851;
assign addr[24017]= 1743623590;
assign addr[24018]= 1787159411;
assign addr[24019]= 1828428082;
assign addr[24020]= 1867377253;
assign addr[24021]= 1903957513;
assign addr[24022]= 1938122457;
assign addr[24023]= 1969828744;
assign addr[24024]= 1999036154;
assign addr[24025]= 2025707632;
assign addr[24026]= 2049809346;
assign addr[24027]= 2071310720;
assign addr[24028]= 2090184478;
assign addr[24029]= 2106406677;
assign addr[24030]= 2119956737;
assign addr[24031]= 2130817471;
assign addr[24032]= 2138975100;
assign addr[24033]= 2144419275;
assign addr[24034]= 2147143090;
assign addr[24035]= 2147143090;
assign addr[24036]= 2144419275;
assign addr[24037]= 2138975100;
assign addr[24038]= 2130817471;
assign addr[24039]= 2119956737;
assign addr[24040]= 2106406677;
assign addr[24041]= 2090184478;
assign addr[24042]= 2071310720;
assign addr[24043]= 2049809346;
assign addr[24044]= 2025707632;
assign addr[24045]= 1999036154;
assign addr[24046]= 1969828744;
assign addr[24047]= 1938122457;
assign addr[24048]= 1903957513;
assign addr[24049]= 1867377253;
assign addr[24050]= 1828428082;
assign addr[24051]= 1787159411;
assign addr[24052]= 1743623590;
assign addr[24053]= 1697875851;
assign addr[24054]= 1649974225;
assign addr[24055]= 1599979481;
assign addr[24056]= 1547955041;
assign addr[24057]= 1493966902;
assign addr[24058]= 1438083551;
assign addr[24059]= 1380375881;
assign addr[24060]= 1320917099;
assign addr[24061]= 1259782632;
assign addr[24062]= 1197050035;
assign addr[24063]= 1132798888;
assign addr[24064]= 1067110699;
assign addr[24065]= 1000068799;
assign addr[24066]= 931758235;
assign addr[24067]= 862265664;
assign addr[24068]= 791679244;
assign addr[24069]= 720088517;
assign addr[24070]= 647584304;
assign addr[24071]= 574258580;
assign addr[24072]= 500204365;
assign addr[24073]= 425515602;
assign addr[24074]= 350287041;
assign addr[24075]= 274614114;
assign addr[24076]= 198592817;
assign addr[24077]= 122319591;
assign addr[24078]= 45891193;
assign addr[24079]= -30595422;
assign addr[24080]= -107043224;
assign addr[24081]= -183355234;
assign addr[24082]= -259434643;
assign addr[24083]= -335184940;
assign addr[24084]= -410510029;
assign addr[24085]= -485314355;
assign addr[24086]= -559503022;
assign addr[24087]= -632981917;
assign addr[24088]= -705657826;
assign addr[24089]= -777438554;
assign addr[24090]= -848233042;
assign addr[24091]= -917951481;
assign addr[24092]= -986505429;
assign addr[24093]= -1053807919;
assign addr[24094]= -1119773573;
assign addr[24095]= -1184318708;
assign addr[24096]= -1247361445;
assign addr[24097]= -1308821808;
assign addr[24098]= -1368621831;
assign addr[24099]= -1426685652;
assign addr[24100]= -1482939614;
assign addr[24101]= -1537312353;
assign addr[24102]= -1589734894;
assign addr[24103]= -1640140734;
assign addr[24104]= -1688465931;
assign addr[24105]= -1734649179;
assign addr[24106]= -1778631892;
assign addr[24107]= -1820358275;
assign addr[24108]= -1859775393;
assign addr[24109]= -1896833245;
assign addr[24110]= -1931484818;
assign addr[24111]= -1963686155;
assign addr[24112]= -1993396407;
assign addr[24113]= -2020577882;
assign addr[24114]= -2045196100;
assign addr[24115]= -2067219829;
assign addr[24116]= -2086621133;
assign addr[24117]= -2103375398;
assign addr[24118]= -2117461370;
assign addr[24119]= -2128861181;
assign addr[24120]= -2137560369;
assign addr[24121]= -2143547897;
assign addr[24122]= -2146816171;
assign addr[24123]= -2147361045;
assign addr[24124]= -2145181827;
assign addr[24125]= -2140281282;
assign addr[24126]= -2132665626;
assign addr[24127]= -2122344521;
assign addr[24128]= -2109331059;
assign addr[24129]= -2093641749;
assign addr[24130]= -2075296495;
assign addr[24131]= -2054318569;
assign addr[24132]= -2030734582;
assign addr[24133]= -2004574453;
assign addr[24134]= -1975871368;
assign addr[24135]= -1944661739;
assign addr[24136]= -1910985158;
assign addr[24137]= -1874884346;
assign addr[24138]= -1836405100;
assign addr[24139]= -1795596234;
assign addr[24140]= -1752509516;
assign addr[24141]= -1707199606;
assign addr[24142]= -1659723983;
assign addr[24143]= -1610142873;
assign addr[24144]= -1558519173;
assign addr[24145]= -1504918373;
assign addr[24146]= -1449408469;
assign addr[24147]= -1392059879;
assign addr[24148]= -1332945355;
assign addr[24149]= -1272139887;
assign addr[24150]= -1209720613;
assign addr[24151]= -1145766716;
assign addr[24152]= -1080359326;
assign addr[24153]= -1013581418;
assign addr[24154]= -945517704;
assign addr[24155]= -876254528;
assign addr[24156]= -805879757;
assign addr[24157]= -734482665;
assign addr[24158]= -662153826;
assign addr[24159]= -588984994;
assign addr[24160]= -515068990;
assign addr[24161]= -440499581;
assign addr[24162]= -365371365;
assign addr[24163]= -289779648;
assign addr[24164]= -213820322;
assign addr[24165]= -137589750;
assign addr[24166]= -61184634;
assign addr[24167]= 15298099;
assign addr[24168]= 91761426;
assign addr[24169]= 168108346;
assign addr[24170]= 244242007;
assign addr[24171]= 320065829;
assign addr[24172]= 395483624;
assign addr[24173]= 470399716;
assign addr[24174]= 544719071;
assign addr[24175]= 618347408;
assign addr[24176]= 691191324;
assign addr[24177]= 763158411;
assign addr[24178]= 834157373;
assign addr[24179]= 904098143;
assign addr[24180]= 972891995;
assign addr[24181]= 1040451659;
assign addr[24182]= 1106691431;
assign addr[24183]= 1171527280;
assign addr[24184]= 1234876957;
assign addr[24185]= 1296660098;
assign addr[24186]= 1356798326;
assign addr[24187]= 1415215352;
assign addr[24188]= 1471837070;
assign addr[24189]= 1526591649;
assign addr[24190]= 1579409630;
assign addr[24191]= 1630224009;
assign addr[24192]= 1678970324;
assign addr[24193]= 1725586737;
assign addr[24194]= 1770014111;
assign addr[24195]= 1812196087;
assign addr[24196]= 1852079154;
assign addr[24197]= 1889612716;
assign addr[24198]= 1924749160;
assign addr[24199]= 1957443913;
assign addr[24200]= 1987655498;
assign addr[24201]= 2015345591;
assign addr[24202]= 2040479063;
assign addr[24203]= 2063024031;
assign addr[24204]= 2082951896;
assign addr[24205]= 2100237377;
assign addr[24206]= 2114858546;
assign addr[24207]= 2126796855;
assign addr[24208]= 2136037160;
assign addr[24209]= 2142567738;
assign addr[24210]= 2146380306;
assign addr[24211]= 2147470025;
assign addr[24212]= 2145835515;
assign addr[24213]= 2141478848;
assign addr[24214]= 2134405552;
assign addr[24215]= 2124624598;
assign addr[24216]= 2112148396;
assign addr[24217]= 2096992772;
assign addr[24218]= 2079176953;
assign addr[24219]= 2058723538;
assign addr[24220]= 2035658475;
assign addr[24221]= 2010011024;
assign addr[24222]= 1981813720;
assign addr[24223]= 1951102334;
assign addr[24224]= 1917915825;
assign addr[24225]= 1882296293;
assign addr[24226]= 1844288924;
assign addr[24227]= 1803941934;
assign addr[24228]= 1761306505;
assign addr[24229]= 1716436725;
assign addr[24230]= 1669389513;
assign addr[24231]= 1620224553;
assign addr[24232]= 1569004214;
assign addr[24233]= 1515793473;
assign addr[24234]= 1460659832;
assign addr[24235]= 1403673233;
assign addr[24236]= 1344905966;
assign addr[24237]= 1284432584;
assign addr[24238]= 1222329801;
assign addr[24239]= 1158676398;
assign addr[24240]= 1093553126;
assign addr[24241]= 1027042599;
assign addr[24242]= 959229189;
assign addr[24243]= 890198924;
assign addr[24244]= 820039373;
assign addr[24245]= 748839539;
assign addr[24246]= 676689746;
assign addr[24247]= 603681519;
assign addr[24248]= 529907477;
assign addr[24249]= 455461206;
assign addr[24250]= 380437148;
assign addr[24251]= 304930476;
assign addr[24252]= 229036977;
assign addr[24253]= 152852926;
assign addr[24254]= 76474970;
assign addr[24255]= 0;
assign addr[24256]= -76474970;
assign addr[24257]= -152852926;
assign addr[24258]= -229036977;
assign addr[24259]= -304930476;
assign addr[24260]= -380437148;
assign addr[24261]= -455461206;
assign addr[24262]= -529907477;
assign addr[24263]= -603681519;
assign addr[24264]= -676689746;
assign addr[24265]= -748839539;
assign addr[24266]= -820039373;
assign addr[24267]= -890198924;
assign addr[24268]= -959229189;
assign addr[24269]= -1027042599;
assign addr[24270]= -1093553126;
assign addr[24271]= -1158676398;
assign addr[24272]= -1222329801;
assign addr[24273]= -1284432584;
assign addr[24274]= -1344905966;
assign addr[24275]= -1403673233;
assign addr[24276]= -1460659832;
assign addr[24277]= -1515793473;
assign addr[24278]= -1569004214;
assign addr[24279]= -1620224553;
assign addr[24280]= -1669389513;
assign addr[24281]= -1716436725;
assign addr[24282]= -1761306505;
assign addr[24283]= -1803941934;
assign addr[24284]= -1844288924;
assign addr[24285]= -1882296293;
assign addr[24286]= -1917915825;
assign addr[24287]= -1951102334;
assign addr[24288]= -1981813720;
assign addr[24289]= -2010011024;
assign addr[24290]= -2035658475;
assign addr[24291]= -2058723538;
assign addr[24292]= -2079176953;
assign addr[24293]= -2096992772;
assign addr[24294]= -2112148396;
assign addr[24295]= -2124624598;
assign addr[24296]= -2134405552;
assign addr[24297]= -2141478848;
assign addr[24298]= -2145835515;
assign addr[24299]= -2147470025;
assign addr[24300]= -2146380306;
assign addr[24301]= -2142567738;
assign addr[24302]= -2136037160;
assign addr[24303]= -2126796855;
assign addr[24304]= -2114858546;
assign addr[24305]= -2100237377;
assign addr[24306]= -2082951896;
assign addr[24307]= -2063024031;
assign addr[24308]= -2040479063;
assign addr[24309]= -2015345591;
assign addr[24310]= -1987655498;
assign addr[24311]= -1957443913;
assign addr[24312]= -1924749160;
assign addr[24313]= -1889612716;
assign addr[24314]= -1852079154;
assign addr[24315]= -1812196087;
assign addr[24316]= -1770014111;
assign addr[24317]= -1725586737;
assign addr[24318]= -1678970324;
assign addr[24319]= -1630224009;
assign addr[24320]= -1579409630;
assign addr[24321]= -1526591649;
assign addr[24322]= -1471837070;
assign addr[24323]= -1415215352;
assign addr[24324]= -1356798326;
assign addr[24325]= -1296660098;
assign addr[24326]= -1234876957;
assign addr[24327]= -1171527280;
assign addr[24328]= -1106691431;
assign addr[24329]= -1040451659;
assign addr[24330]= -972891995;
assign addr[24331]= -904098143;
assign addr[24332]= -834157373;
assign addr[24333]= -763158411;
assign addr[24334]= -691191324;
assign addr[24335]= -618347408;
assign addr[24336]= -544719071;
assign addr[24337]= -470399716;
assign addr[24338]= -395483624;
assign addr[24339]= -320065829;
assign addr[24340]= -244242007;
assign addr[24341]= -168108346;
assign addr[24342]= -91761426;
assign addr[24343]= -15298099;
assign addr[24344]= 61184634;
assign addr[24345]= 137589750;
assign addr[24346]= 213820322;
assign addr[24347]= 289779648;
assign addr[24348]= 365371365;
assign addr[24349]= 440499581;
assign addr[24350]= 515068990;
assign addr[24351]= 588984994;
assign addr[24352]= 662153826;
assign addr[24353]= 734482665;
assign addr[24354]= 805879757;
assign addr[24355]= 876254528;
assign addr[24356]= 945517704;
assign addr[24357]= 1013581418;
assign addr[24358]= 1080359326;
assign addr[24359]= 1145766716;
assign addr[24360]= 1209720613;
assign addr[24361]= 1272139887;
assign addr[24362]= 1332945355;
assign addr[24363]= 1392059879;
assign addr[24364]= 1449408469;
assign addr[24365]= 1504918373;
assign addr[24366]= 1558519173;
assign addr[24367]= 1610142873;
assign addr[24368]= 1659723983;
assign addr[24369]= 1707199606;
assign addr[24370]= 1752509516;
assign addr[24371]= 1795596234;
assign addr[24372]= 1836405100;
assign addr[24373]= 1874884346;
assign addr[24374]= 1910985158;
assign addr[24375]= 1944661739;
assign addr[24376]= 1975871368;
assign addr[24377]= 2004574453;
assign addr[24378]= 2030734582;
assign addr[24379]= 2054318569;
assign addr[24380]= 2075296495;
assign addr[24381]= 2093641749;
assign addr[24382]= 2109331059;
assign addr[24383]= 2122344521;
assign addr[24384]= 2132665626;
assign addr[24385]= 2140281282;
assign addr[24386]= 2145181827;
assign addr[24387]= 2147361045;
assign addr[24388]= 2146816171;
assign addr[24389]= 2143547897;
assign addr[24390]= 2137560369;
assign addr[24391]= 2128861181;
assign addr[24392]= 2117461370;
assign addr[24393]= 2103375398;
assign addr[24394]= 2086621133;
assign addr[24395]= 2067219829;
assign addr[24396]= 2045196100;
assign addr[24397]= 2020577882;
assign addr[24398]= 1993396407;
assign addr[24399]= 1963686155;
assign addr[24400]= 1931484818;
assign addr[24401]= 1896833245;
assign addr[24402]= 1859775393;
assign addr[24403]= 1820358275;
assign addr[24404]= 1778631892;
assign addr[24405]= 1734649179;
assign addr[24406]= 1688465931;
assign addr[24407]= 1640140734;
assign addr[24408]= 1589734894;
assign addr[24409]= 1537312353;
assign addr[24410]= 1482939614;
assign addr[24411]= 1426685652;
assign addr[24412]= 1368621831;
assign addr[24413]= 1308821808;
assign addr[24414]= 1247361445;
assign addr[24415]= 1184318708;
assign addr[24416]= 1119773573;
assign addr[24417]= 1053807919;
assign addr[24418]= 986505429;
assign addr[24419]= 917951481;
assign addr[24420]= 848233042;
assign addr[24421]= 777438554;
assign addr[24422]= 705657826;
assign addr[24423]= 632981917;
assign addr[24424]= 559503022;
assign addr[24425]= 485314355;
assign addr[24426]= 410510029;
assign addr[24427]= 335184940;
assign addr[24428]= 259434643;
assign addr[24429]= 183355234;
assign addr[24430]= 107043224;
assign addr[24431]= 30595422;
assign addr[24432]= -45891193;
assign addr[24433]= -122319591;
assign addr[24434]= -198592817;
assign addr[24435]= -274614114;
assign addr[24436]= -350287041;
assign addr[24437]= -425515602;
assign addr[24438]= -500204365;
assign addr[24439]= -574258580;
assign addr[24440]= -647584304;
assign addr[24441]= -720088517;
assign addr[24442]= -791679244;
assign addr[24443]= -862265664;
assign addr[24444]= -931758235;
assign addr[24445]= -1000068799;
assign addr[24446]= -1067110699;
assign addr[24447]= -1132798888;
assign addr[24448]= -1197050035;
assign addr[24449]= -1259782632;
assign addr[24450]= -1320917099;
assign addr[24451]= -1380375881;
assign addr[24452]= -1438083551;
assign addr[24453]= -1493966902;
assign addr[24454]= -1547955041;
assign addr[24455]= -1599979481;
assign addr[24456]= -1649974225;
assign addr[24457]= -1697875851;
assign addr[24458]= -1743623590;
assign addr[24459]= -1787159411;
assign addr[24460]= -1828428082;
assign addr[24461]= -1867377253;
assign addr[24462]= -1903957513;
assign addr[24463]= -1938122457;
assign addr[24464]= -1969828744;
assign addr[24465]= -1999036154;
assign addr[24466]= -2025707632;
assign addr[24467]= -2049809346;
assign addr[24468]= -2071310720;
assign addr[24469]= -2090184478;
assign addr[24470]= -2106406677;
assign addr[24471]= -2119956737;
assign addr[24472]= -2130817471;
assign addr[24473]= -2138975100;
assign addr[24474]= -2144419275;
assign addr[24475]= -2147143090;
assign addr[24476]= -2147143090;
assign addr[24477]= -2144419275;
assign addr[24478]= -2138975100;
assign addr[24479]= -2130817471;
assign addr[24480]= -2119956737;
assign addr[24481]= -2106406677;
assign addr[24482]= -2090184478;
assign addr[24483]= -2071310720;
assign addr[24484]= -2049809346;
assign addr[24485]= -2025707632;
assign addr[24486]= -1999036154;
assign addr[24487]= -1969828744;
assign addr[24488]= -1938122457;
assign addr[24489]= -1903957513;
assign addr[24490]= -1867377253;
assign addr[24491]= -1828428082;
assign addr[24492]= -1787159411;
assign addr[24493]= -1743623590;
assign addr[24494]= -1697875851;
assign addr[24495]= -1649974225;
assign addr[24496]= -1599979481;
assign addr[24497]= -1547955041;
assign addr[24498]= -1493966902;
assign addr[24499]= -1438083551;
assign addr[24500]= -1380375881;
assign addr[24501]= -1320917099;
assign addr[24502]= -1259782632;
assign addr[24503]= -1197050035;
assign addr[24504]= -1132798888;
assign addr[24505]= -1067110699;
assign addr[24506]= -1000068799;
assign addr[24507]= -931758235;
assign addr[24508]= -862265664;
assign addr[24509]= -791679244;
assign addr[24510]= -720088517;
assign addr[24511]= -647584304;
assign addr[24512]= -574258580;
assign addr[24513]= -500204365;
assign addr[24514]= -425515602;
assign addr[24515]= -350287041;
assign addr[24516]= -274614114;
assign addr[24517]= -198592817;
assign addr[24518]= -122319591;
assign addr[24519]= -45891193;
assign addr[24520]= 30595422;
assign addr[24521]= 107043224;
assign addr[24522]= 183355234;
assign addr[24523]= 259434643;
assign addr[24524]= 335184940;
assign addr[24525]= 410510029;
assign addr[24526]= 485314355;
assign addr[24527]= 559503022;
assign addr[24528]= 632981917;
assign addr[24529]= 705657826;
assign addr[24530]= 777438554;
assign addr[24531]= 848233042;
assign addr[24532]= 917951481;
assign addr[24533]= 986505429;
assign addr[24534]= 1053807919;
assign addr[24535]= 1119773573;
assign addr[24536]= 1184318708;
assign addr[24537]= 1247361445;
assign addr[24538]= 1308821808;
assign addr[24539]= 1368621831;
assign addr[24540]= 1426685652;
assign addr[24541]= 1482939614;
assign addr[24542]= 1537312353;
assign addr[24543]= 1589734894;
assign addr[24544]= 1640140734;
assign addr[24545]= 1688465931;
assign addr[24546]= 1734649179;
assign addr[24547]= 1778631892;
assign addr[24548]= 1820358275;
assign addr[24549]= 1859775393;
assign addr[24550]= 1896833245;
assign addr[24551]= 1931484818;
assign addr[24552]= 1963686155;
assign addr[24553]= 1993396407;
assign addr[24554]= 2020577882;
assign addr[24555]= 2045196100;
assign addr[24556]= 2067219829;
assign addr[24557]= 2086621133;
assign addr[24558]= 2103375398;
assign addr[24559]= 2117461370;
assign addr[24560]= 2128861181;
assign addr[24561]= 2137560369;
assign addr[24562]= 2143547897;
assign addr[24563]= 2146816171;
assign addr[24564]= 2147361045;
assign addr[24565]= 2145181827;
assign addr[24566]= 2140281282;
assign addr[24567]= 2132665626;
assign addr[24568]= 2122344521;
assign addr[24569]= 2109331059;
assign addr[24570]= 2093641749;
assign addr[24571]= 2075296495;
assign addr[24572]= 2054318569;
assign addr[24573]= 2030734582;
assign addr[24574]= 2004574453;
assign addr[24575]= 1975871368;
assign addr[24576]= 1944661739;
assign addr[24577]= 1910985158;
assign addr[24578]= 1874884346;
assign addr[24579]= 1836405100;
assign addr[24580]= 1795596234;
assign addr[24581]= 1752509516;
assign addr[24582]= 1707199606;
assign addr[24583]= 1659723983;
assign addr[24584]= 1610142873;
assign addr[24585]= 1558519173;
assign addr[24586]= 1504918373;
assign addr[24587]= 1449408469;
assign addr[24588]= 1392059879;
assign addr[24589]= 1332945355;
assign addr[24590]= 1272139887;
assign addr[24591]= 1209720613;
assign addr[24592]= 1145766716;
assign addr[24593]= 1080359326;
assign addr[24594]= 1013581418;
assign addr[24595]= 945517704;
assign addr[24596]= 876254528;
assign addr[24597]= 805879757;
assign addr[24598]= 734482665;
assign addr[24599]= 662153826;
assign addr[24600]= 588984994;
assign addr[24601]= 515068990;
assign addr[24602]= 440499581;
assign addr[24603]= 365371365;
assign addr[24604]= 289779648;
assign addr[24605]= 213820322;
assign addr[24606]= 137589750;
assign addr[24607]= 61184634;
assign addr[24608]= -15298099;
assign addr[24609]= -91761426;
assign addr[24610]= -168108346;
assign addr[24611]= -244242007;
assign addr[24612]= -320065829;
assign addr[24613]= -395483624;
assign addr[24614]= -470399716;
assign addr[24615]= -544719071;
assign addr[24616]= -618347408;
assign addr[24617]= -691191324;
assign addr[24618]= -763158411;
assign addr[24619]= -834157373;
assign addr[24620]= -904098143;
assign addr[24621]= -972891995;
assign addr[24622]= -1040451659;
assign addr[24623]= -1106691431;
assign addr[24624]= -1171527280;
assign addr[24625]= -1234876957;
assign addr[24626]= -1296660098;
assign addr[24627]= -1356798326;
assign addr[24628]= -1415215352;
assign addr[24629]= -1471837070;
assign addr[24630]= -1526591649;
assign addr[24631]= -1579409630;
assign addr[24632]= -1630224009;
assign addr[24633]= -1678970324;
assign addr[24634]= -1725586737;
assign addr[24635]= -1770014111;
assign addr[24636]= -1812196087;
assign addr[24637]= -1852079154;
assign addr[24638]= -1889612716;
assign addr[24639]= -1924749160;
assign addr[24640]= -1957443913;
assign addr[24641]= -1987655498;
assign addr[24642]= -2015345591;
assign addr[24643]= -2040479063;
assign addr[24644]= -2063024031;
assign addr[24645]= -2082951896;
assign addr[24646]= -2100237377;
assign addr[24647]= -2114858546;
assign addr[24648]= -2126796855;
assign addr[24649]= -2136037160;
assign addr[24650]= -2142567738;
assign addr[24651]= -2146380306;
assign addr[24652]= -2147470025;
assign addr[24653]= -2145835515;
assign addr[24654]= -2141478848;
assign addr[24655]= -2134405552;
assign addr[24656]= -2124624598;
assign addr[24657]= -2112148396;
assign addr[24658]= -2096992772;
assign addr[24659]= -2079176953;
assign addr[24660]= -2058723538;
assign addr[24661]= -2035658475;
assign addr[24662]= -2010011024;
assign addr[24663]= -1981813720;
assign addr[24664]= -1951102334;
assign addr[24665]= -1917915825;
assign addr[24666]= -1882296293;
assign addr[24667]= -1844288924;
assign addr[24668]= -1803941934;
assign addr[24669]= -1761306505;
assign addr[24670]= -1716436725;
assign addr[24671]= -1669389513;
assign addr[24672]= -1620224553;
assign addr[24673]= -1569004214;
assign addr[24674]= -1515793473;
assign addr[24675]= -1460659832;
assign addr[24676]= -1403673233;
assign addr[24677]= -1344905966;
assign addr[24678]= -1284432584;
assign addr[24679]= -1222329801;
assign addr[24680]= -1158676398;
assign addr[24681]= -1093553126;
assign addr[24682]= -1027042599;
assign addr[24683]= -959229189;
assign addr[24684]= -890198924;
assign addr[24685]= -820039373;
assign addr[24686]= -748839539;
assign addr[24687]= -676689746;
assign addr[24688]= -603681519;
assign addr[24689]= -529907477;
assign addr[24690]= -455461206;
assign addr[24691]= -380437148;
assign addr[24692]= -304930476;
assign addr[24693]= -229036977;
assign addr[24694]= -152852926;
assign addr[24695]= -76474970;
assign addr[24696]= 0;
assign addr[24697]= 76474970;
assign addr[24698]= 152852926;
assign addr[24699]= 229036977;
assign addr[24700]= 304930476;
assign addr[24701]= 380437148;
assign addr[24702]= 455461206;
assign addr[24703]= 529907477;
assign addr[24704]= 603681519;
assign addr[24705]= 676689746;
assign addr[24706]= 748839539;
assign addr[24707]= 820039373;
assign addr[24708]= 890198924;
assign addr[24709]= 959229189;
assign addr[24710]= 1027042599;
assign addr[24711]= 1093553126;
assign addr[24712]= 1158676398;
assign addr[24713]= 1222329801;
assign addr[24714]= 1284432584;
assign addr[24715]= 1344905966;
assign addr[24716]= 1403673233;
assign addr[24717]= 1460659832;
assign addr[24718]= 1515793473;
assign addr[24719]= 1569004214;
assign addr[24720]= 1620224553;
assign addr[24721]= 1669389513;
assign addr[24722]= 1716436725;
assign addr[24723]= 1761306505;
assign addr[24724]= 1803941934;
assign addr[24725]= 1844288924;
assign addr[24726]= 1882296293;
assign addr[24727]= 1917915825;
assign addr[24728]= 1951102334;
assign addr[24729]= 1981813720;
assign addr[24730]= 2010011024;
assign addr[24731]= 2035658475;
assign addr[24732]= 2058723538;
assign addr[24733]= 2079176953;
assign addr[24734]= 2096992772;
assign addr[24735]= 2112148396;
assign addr[24736]= 2124624598;
assign addr[24737]= 2134405552;
assign addr[24738]= 2141478848;
assign addr[24739]= 2145835515;
assign addr[24740]= 2147470025;
assign addr[24741]= 2146380306;
assign addr[24742]= 2142567738;
assign addr[24743]= 2136037160;
assign addr[24744]= 2126796855;
assign addr[24745]= 2114858546;
assign addr[24746]= 2100237377;
assign addr[24747]= 2082951896;
assign addr[24748]= 2063024031;
assign addr[24749]= 2040479063;
assign addr[24750]= 2015345591;
assign addr[24751]= 1987655498;
assign addr[24752]= 1957443913;
assign addr[24753]= 1924749160;
assign addr[24754]= 1889612716;
assign addr[24755]= 1852079154;
assign addr[24756]= 1812196087;
assign addr[24757]= 1770014111;
assign addr[24758]= 1725586737;
assign addr[24759]= 1678970324;
assign addr[24760]= 1630224009;
assign addr[24761]= 1579409630;
assign addr[24762]= 1526591649;
assign addr[24763]= 1471837070;
assign addr[24764]= 1415215352;
assign addr[24765]= 1356798326;
assign addr[24766]= 1296660098;
assign addr[24767]= 1234876957;
assign addr[24768]= 1171527280;
assign addr[24769]= 1106691431;
assign addr[24770]= 1040451659;
assign addr[24771]= 972891995;
assign addr[24772]= 904098143;
assign addr[24773]= 834157373;
assign addr[24774]= 763158411;
assign addr[24775]= 691191324;
assign addr[24776]= 618347408;
assign addr[24777]= 544719071;
assign addr[24778]= 470399716;
assign addr[24779]= 395483624;
assign addr[24780]= 320065829;
assign addr[24781]= 244242007;
assign addr[24782]= 168108346;
assign addr[24783]= 91761426;
assign addr[24784]= 15298099;
assign addr[24785]= -61184634;
assign addr[24786]= -137589750;
assign addr[24787]= -213820322;
assign addr[24788]= -289779648;
assign addr[24789]= -365371365;
assign addr[24790]= -440499581;
assign addr[24791]= -515068990;
assign addr[24792]= -588984994;
assign addr[24793]= -662153826;
assign addr[24794]= -734482665;
assign addr[24795]= -805879757;
assign addr[24796]= -876254528;
assign addr[24797]= -945517704;
assign addr[24798]= -1013581418;
assign addr[24799]= -1080359326;
assign addr[24800]= -1145766716;
assign addr[24801]= -1209720613;
assign addr[24802]= -1272139887;
assign addr[24803]= -1332945355;
assign addr[24804]= -1392059879;
assign addr[24805]= -1449408469;
assign addr[24806]= -1504918373;
assign addr[24807]= -1558519173;
assign addr[24808]= -1610142873;
assign addr[24809]= -1659723983;
assign addr[24810]= -1707199606;
assign addr[24811]= -1752509516;
assign addr[24812]= -1795596234;
assign addr[24813]= -1836405100;
assign addr[24814]= -1874884346;
assign addr[24815]= -1910985158;
assign addr[24816]= -1944661739;
assign addr[24817]= -1975871368;
assign addr[24818]= -2004574453;
assign addr[24819]= -2030734582;
assign addr[24820]= -2054318569;
assign addr[24821]= -2075296495;
assign addr[24822]= -2093641749;
assign addr[24823]= -2109331059;
assign addr[24824]= -2122344521;
assign addr[24825]= -2132665626;
assign addr[24826]= -2140281282;
assign addr[24827]= -2145181827;
assign addr[24828]= -2147361045;
assign addr[24829]= -2146816171;
assign addr[24830]= -2143547897;
assign addr[24831]= -2137560369;
assign addr[24832]= -2128861181;
assign addr[24833]= -2117461370;
assign addr[24834]= -2103375398;
assign addr[24835]= -2086621133;
assign addr[24836]= -2067219829;
assign addr[24837]= -2045196100;
assign addr[24838]= -2020577882;
assign addr[24839]= -1993396407;
assign addr[24840]= -1963686155;
assign addr[24841]= -1931484818;
assign addr[24842]= -1896833245;
assign addr[24843]= -1859775393;
assign addr[24844]= -1820358275;
assign addr[24845]= -1778631892;
assign addr[24846]= -1734649179;
assign addr[24847]= -1688465931;
assign addr[24848]= -1640140734;
assign addr[24849]= -1589734894;
assign addr[24850]= -1537312353;
assign addr[24851]= -1482939614;
assign addr[24852]= -1426685652;
assign addr[24853]= -1368621831;
assign addr[24854]= -1308821808;
assign addr[24855]= -1247361445;
assign addr[24856]= -1184318708;
assign addr[24857]= -1119773573;
assign addr[24858]= -1053807919;
assign addr[24859]= -986505429;
assign addr[24860]= -917951481;
assign addr[24861]= -848233042;
assign addr[24862]= -777438554;
assign addr[24863]= -705657826;
assign addr[24864]= -632981917;
assign addr[24865]= -559503022;
assign addr[24866]= -485314355;
assign addr[24867]= -410510029;
assign addr[24868]= -335184940;
assign addr[24869]= -259434643;
assign addr[24870]= -183355234;
assign addr[24871]= -107043224;
assign addr[24872]= -30595422;
assign addr[24873]= 45891193;
assign addr[24874]= 122319591;
assign addr[24875]= 198592817;
assign addr[24876]= 274614114;
assign addr[24877]= 350287041;
assign addr[24878]= 425515602;
assign addr[24879]= 500204365;
assign addr[24880]= 574258580;
assign addr[24881]= 647584304;
assign addr[24882]= 720088517;
assign addr[24883]= 791679244;
assign addr[24884]= 862265664;
assign addr[24885]= 931758235;
assign addr[24886]= 1000068799;
assign addr[24887]= 1067110699;
assign addr[24888]= 1132798888;
assign addr[24889]= 1197050035;
assign addr[24890]= 1259782632;
assign addr[24891]= 1320917099;
assign addr[24892]= 1380375881;
assign addr[24893]= 1438083551;
assign addr[24894]= 1493966902;
assign addr[24895]= 1547955041;
assign addr[24896]= 1599979481;
assign addr[24897]= 1649974225;
assign addr[24898]= 1697875851;
assign addr[24899]= 1743623590;
assign addr[24900]= 1787159411;
assign addr[24901]= 1828428082;
assign addr[24902]= 1867377253;
assign addr[24903]= 1903957513;
assign addr[24904]= 1938122457;
assign addr[24905]= 1969828744;
assign addr[24906]= 1999036154;
assign addr[24907]= 2025707632;
assign addr[24908]= 2049809346;
assign addr[24909]= 2071310720;
assign addr[24910]= 2090184478;
assign addr[24911]= 2106406677;
assign addr[24912]= 2119956737;
assign addr[24913]= 2130817471;
assign addr[24914]= 2138975100;
assign addr[24915]= 2144419275;
assign addr[24916]= 2147143090;
assign addr[24917]= 2147143090;
assign addr[24918]= 2144419275;
assign addr[24919]= 2138975100;
assign addr[24920]= 2130817471;
assign addr[24921]= 2119956737;
assign addr[24922]= 2106406677;
assign addr[24923]= 2090184478;
assign addr[24924]= 2071310720;
assign addr[24925]= 2049809346;
assign addr[24926]= 2025707632;
assign addr[24927]= 1999036154;
assign addr[24928]= 1969828744;
assign addr[24929]= 1938122457;
assign addr[24930]= 1903957513;
assign addr[24931]= 1867377253;
assign addr[24932]= 1828428082;
assign addr[24933]= 1787159411;
assign addr[24934]= 1743623590;
assign addr[24935]= 1697875851;
assign addr[24936]= 1649974225;
assign addr[24937]= 1599979481;
assign addr[24938]= 1547955041;
assign addr[24939]= 1493966902;
assign addr[24940]= 1438083551;
assign addr[24941]= 1380375881;
assign addr[24942]= 1320917099;
assign addr[24943]= 1259782632;
assign addr[24944]= 1197050035;
assign addr[24945]= 1132798888;
assign addr[24946]= 1067110699;
assign addr[24947]= 1000068799;
assign addr[24948]= 931758235;
assign addr[24949]= 862265664;
assign addr[24950]= 791679244;
assign addr[24951]= 720088517;
assign addr[24952]= 647584304;
assign addr[24953]= 574258580;
assign addr[24954]= 500204365;
assign addr[24955]= 425515602;
assign addr[24956]= 350287041;
assign addr[24957]= 274614114;
assign addr[24958]= 198592817;
assign addr[24959]= 122319591;
assign addr[24960]= 45891193;
assign addr[24961]= -30595422;
assign addr[24962]= -107043224;
assign addr[24963]= -183355234;
assign addr[24964]= -259434643;
assign addr[24965]= -335184940;
assign addr[24966]= -410510029;
assign addr[24967]= -485314355;
assign addr[24968]= -559503022;
assign addr[24969]= -632981917;
assign addr[24970]= -705657826;
assign addr[24971]= -777438554;
assign addr[24972]= -848233042;
assign addr[24973]= -917951481;
assign addr[24974]= -986505429;
assign addr[24975]= -1053807919;
assign addr[24976]= -1119773573;
assign addr[24977]= -1184318708;
assign addr[24978]= -1247361445;
assign addr[24979]= -1308821808;
assign addr[24980]= -1368621831;
assign addr[24981]= -1426685652;
assign addr[24982]= -1482939614;
assign addr[24983]= -1537312353;
assign addr[24984]= -1589734894;
assign addr[24985]= -1640140734;
assign addr[24986]= -1688465931;
assign addr[24987]= -1734649179;
assign addr[24988]= -1778631892;
assign addr[24989]= -1820358275;
assign addr[24990]= -1859775393;
assign addr[24991]= -1896833245;
assign addr[24992]= -1931484818;
assign addr[24993]= -1963686155;
assign addr[24994]= -1993396407;
assign addr[24995]= -2020577882;
assign addr[24996]= -2045196100;
assign addr[24997]= -2067219829;
assign addr[24998]= -2086621133;
assign addr[24999]= -2103375398;
assign addr[25000]= -2117461370;
assign addr[25001]= -2128861181;
assign addr[25002]= -2137560369;
assign addr[25003]= -2143547897;
assign addr[25004]= -2146816171;
assign addr[25005]= -2147361045;
assign addr[25006]= -2145181827;
assign addr[25007]= -2140281282;
assign addr[25008]= -2132665626;
assign addr[25009]= -2122344521;
assign addr[25010]= -2109331059;
assign addr[25011]= -2093641749;
assign addr[25012]= -2075296495;
assign addr[25013]= -2054318569;
assign addr[25014]= -2030734582;
assign addr[25015]= -2004574453;
assign addr[25016]= -1975871368;
assign addr[25017]= -1944661739;
assign addr[25018]= -1910985158;
assign addr[25019]= -1874884346;
assign addr[25020]= -1836405100;
assign addr[25021]= -1795596234;
assign addr[25022]= -1752509516;
assign addr[25023]= -1707199606;
assign addr[25024]= -1659723983;
assign addr[25025]= -1610142873;
assign addr[25026]= -1558519173;
assign addr[25027]= -1504918373;
assign addr[25028]= -1449408469;
assign addr[25029]= -1392059879;
assign addr[25030]= -1332945355;
assign addr[25031]= -1272139887;
assign addr[25032]= -1209720613;
assign addr[25033]= -1145766716;
assign addr[25034]= -1080359326;
assign addr[25035]= -1013581418;
assign addr[25036]= -945517704;
assign addr[25037]= -876254528;
assign addr[25038]= -805879757;
assign addr[25039]= -734482665;
assign addr[25040]= -662153826;
assign addr[25041]= -588984994;
assign addr[25042]= -515068990;
assign addr[25043]= -440499581;
assign addr[25044]= -365371365;
assign addr[25045]= -289779648;
assign addr[25046]= -213820322;
assign addr[25047]= -137589750;
assign addr[25048]= -61184634;
assign addr[25049]= 15298099;
assign addr[25050]= 91761426;
assign addr[25051]= 168108346;
assign addr[25052]= 244242007;
assign addr[25053]= 320065829;
assign addr[25054]= 395483624;
assign addr[25055]= 470399716;
assign addr[25056]= 544719071;
assign addr[25057]= 618347408;
assign addr[25058]= 691191324;
assign addr[25059]= 763158411;
assign addr[25060]= 834157373;
assign addr[25061]= 904098143;
assign addr[25062]= 972891995;
assign addr[25063]= 1040451659;
assign addr[25064]= 1106691431;
assign addr[25065]= 1171527280;
assign addr[25066]= 1234876957;
assign addr[25067]= 1296660098;
assign addr[25068]= 1356798326;
assign addr[25069]= 1415215352;
assign addr[25070]= 1471837070;
assign addr[25071]= 1526591649;
assign addr[25072]= 1579409630;
assign addr[25073]= 1630224009;
assign addr[25074]= 1678970324;
assign addr[25075]= 1725586737;
assign addr[25076]= 1770014111;
assign addr[25077]= 1812196087;
assign addr[25078]= 1852079154;
assign addr[25079]= 1889612716;
assign addr[25080]= 1924749160;
assign addr[25081]= 1957443913;
assign addr[25082]= 1987655498;
assign addr[25083]= 2015345591;
assign addr[25084]= 2040479063;
assign addr[25085]= 2063024031;
assign addr[25086]= 2082951896;
assign addr[25087]= 2100237377;
assign addr[25088]= 2114858546;
assign addr[25089]= 2126796855;
assign addr[25090]= 2136037160;
assign addr[25091]= 2142567738;
assign addr[25092]= 2146380306;
assign addr[25093]= 2147470025;
assign addr[25094]= 2145835515;
assign addr[25095]= 2141478848;
assign addr[25096]= 2134405552;
assign addr[25097]= 2124624598;
assign addr[25098]= 2112148396;
assign addr[25099]= 2096992772;
assign addr[25100]= 2079176953;
assign addr[25101]= 2058723538;
assign addr[25102]= 2035658475;
assign addr[25103]= 2010011024;
assign addr[25104]= 1981813720;
assign addr[25105]= 1951102334;
assign addr[25106]= 1917915825;
assign addr[25107]= 1882296293;
assign addr[25108]= 1844288924;
assign addr[25109]= 1803941934;
assign addr[25110]= 1761306505;
assign addr[25111]= 1716436725;
assign addr[25112]= 1669389513;
assign addr[25113]= 1620224553;
assign addr[25114]= 1569004214;
assign addr[25115]= 1515793473;
assign addr[25116]= 1460659832;
assign addr[25117]= 1403673233;
assign addr[25118]= 1344905966;
assign addr[25119]= 1284432584;
assign addr[25120]= 1222329801;
assign addr[25121]= 1158676398;
assign addr[25122]= 1093553126;
assign addr[25123]= 1027042599;
assign addr[25124]= 959229189;
assign addr[25125]= 890198924;
assign addr[25126]= 820039373;
assign addr[25127]= 748839539;
assign addr[25128]= 676689746;
assign addr[25129]= 603681519;
assign addr[25130]= 529907477;
assign addr[25131]= 455461206;
assign addr[25132]= 380437148;
assign addr[25133]= 304930476;
assign addr[25134]= 229036977;
assign addr[25135]= 152852926;
assign addr[25136]= 76474970;
assign addr[25137]= 0;
assign addr[25138]= -76474970;
assign addr[25139]= -152852926;
assign addr[25140]= -229036977;
assign addr[25141]= -304930476;
assign addr[25142]= -380437148;
assign addr[25143]= -455461206;
assign addr[25144]= -529907477;
assign addr[25145]= -603681519;
assign addr[25146]= -676689746;
assign addr[25147]= -748839539;
assign addr[25148]= -820039373;
assign addr[25149]= -890198924;
assign addr[25150]= -959229189;
assign addr[25151]= -1027042599;
assign addr[25152]= -1093553126;
assign addr[25153]= -1158676398;
assign addr[25154]= -1222329801;
assign addr[25155]= -1284432584;
assign addr[25156]= -1344905966;
assign addr[25157]= -1403673233;
assign addr[25158]= -1460659832;
assign addr[25159]= -1515793473;
assign addr[25160]= -1569004214;
assign addr[25161]= -1620224553;
assign addr[25162]= -1669389513;
assign addr[25163]= -1716436725;
assign addr[25164]= -1761306505;
assign addr[25165]= -1803941934;
assign addr[25166]= -1844288924;
assign addr[25167]= -1882296293;
assign addr[25168]= -1917915825;
assign addr[25169]= -1951102334;
assign addr[25170]= -1981813720;
assign addr[25171]= -2010011024;
assign addr[25172]= -2035658475;
assign addr[25173]= -2058723538;
assign addr[25174]= -2079176953;
assign addr[25175]= -2096992772;
assign addr[25176]= -2112148396;
assign addr[25177]= -2124624598;
assign addr[25178]= -2134405552;
assign addr[25179]= -2141478848;
assign addr[25180]= -2145835515;
assign addr[25181]= -2147470025;
assign addr[25182]= -2146380306;
assign addr[25183]= -2142567738;
assign addr[25184]= -2136037160;
assign addr[25185]= -2126796855;
assign addr[25186]= -2114858546;
assign addr[25187]= -2100237377;
assign addr[25188]= -2082951896;
assign addr[25189]= -2063024031;
assign addr[25190]= -2040479063;
assign addr[25191]= -2015345591;
assign addr[25192]= -1987655498;
assign addr[25193]= -1957443913;
assign addr[25194]= -1924749160;
assign addr[25195]= -1889612716;
assign addr[25196]= -1852079154;
assign addr[25197]= -1812196087;
assign addr[25198]= -1770014111;
assign addr[25199]= -1725586737;
assign addr[25200]= -1678970324;
assign addr[25201]= -1630224009;
assign addr[25202]= -1579409630;
assign addr[25203]= -1526591649;
assign addr[25204]= -1471837070;
assign addr[25205]= -1415215352;
assign addr[25206]= -1356798326;
assign addr[25207]= -1296660098;
assign addr[25208]= -1234876957;
assign addr[25209]= -1171527280;
assign addr[25210]= -1106691431;
assign addr[25211]= -1040451659;
assign addr[25212]= -972891995;
assign addr[25213]= -904098143;
assign addr[25214]= -834157373;
assign addr[25215]= -763158411;
assign addr[25216]= -691191324;
assign addr[25217]= -618347408;
assign addr[25218]= -544719071;
assign addr[25219]= -470399716;
assign addr[25220]= -395483624;
assign addr[25221]= -320065829;
assign addr[25222]= -244242007;
assign addr[25223]= -168108346;
assign addr[25224]= -91761426;
assign addr[25225]= -15298099;
assign addr[25226]= 61184634;
assign addr[25227]= 137589750;
assign addr[25228]= 213820322;
assign addr[25229]= 289779648;
assign addr[25230]= 365371365;
assign addr[25231]= 440499581;
assign addr[25232]= 515068990;
assign addr[25233]= 588984994;
assign addr[25234]= 662153826;
assign addr[25235]= 734482665;
assign addr[25236]= 805879757;
assign addr[25237]= 876254528;
assign addr[25238]= 945517704;
assign addr[25239]= 1013581418;
assign addr[25240]= 1080359326;
assign addr[25241]= 1145766716;
assign addr[25242]= 1209720613;
assign addr[25243]= 1272139887;
assign addr[25244]= 1332945355;
assign addr[25245]= 1392059879;
assign addr[25246]= 1449408469;
assign addr[25247]= 1504918373;
assign addr[25248]= 1558519173;
assign addr[25249]= 1610142873;
assign addr[25250]= 1659723983;
assign addr[25251]= 1707199606;
assign addr[25252]= 1752509516;
assign addr[25253]= 1795596234;
assign addr[25254]= 1836405100;
assign addr[25255]= 1874884346;
assign addr[25256]= 1910985158;
assign addr[25257]= 1944661739;
assign addr[25258]= 1975871368;
assign addr[25259]= 2004574453;
assign addr[25260]= 2030734582;
assign addr[25261]= 2054318569;
assign addr[25262]= 2075296495;
assign addr[25263]= 2093641749;
assign addr[25264]= 2109331059;
assign addr[25265]= 2122344521;
assign addr[25266]= 2132665626;
assign addr[25267]= 2140281282;
assign addr[25268]= 2145181827;
assign addr[25269]= 2147361045;
assign addr[25270]= 2146816171;
assign addr[25271]= 2143547897;
assign addr[25272]= 2137560369;
assign addr[25273]= 2128861181;
assign addr[25274]= 2117461370;
assign addr[25275]= 2103375398;
assign addr[25276]= 2086621133;
assign addr[25277]= 2067219829;
assign addr[25278]= 2045196100;
assign addr[25279]= 2020577882;
assign addr[25280]= 1993396407;
assign addr[25281]= 1963686155;
assign addr[25282]= 1931484818;
assign addr[25283]= 1896833245;
assign addr[25284]= 1859775393;
assign addr[25285]= 1820358275;
assign addr[25286]= 1778631892;
assign addr[25287]= 1734649179;
assign addr[25288]= 1688465931;
assign addr[25289]= 1640140734;
assign addr[25290]= 1589734894;
assign addr[25291]= 1537312353;
assign addr[25292]= 1482939614;
assign addr[25293]= 1426685652;
assign addr[25294]= 1368621831;
assign addr[25295]= 1308821808;
assign addr[25296]= 1247361445;
assign addr[25297]= 1184318708;
assign addr[25298]= 1119773573;
assign addr[25299]= 1053807919;
assign addr[25300]= 986505429;
assign addr[25301]= 917951481;
assign addr[25302]= 848233042;
assign addr[25303]= 777438554;
assign addr[25304]= 705657826;
assign addr[25305]= 632981917;
assign addr[25306]= 559503022;
assign addr[25307]= 485314355;
assign addr[25308]= 410510029;
assign addr[25309]= 335184940;
assign addr[25310]= 259434643;
assign addr[25311]= 183355234;
assign addr[25312]= 107043224;
assign addr[25313]= 30595422;
assign addr[25314]= -45891193;
assign addr[25315]= -122319591;
assign addr[25316]= -198592817;
assign addr[25317]= -274614114;
assign addr[25318]= -350287041;
assign addr[25319]= -425515602;
assign addr[25320]= -500204365;
assign addr[25321]= -574258580;
assign addr[25322]= -647584304;
assign addr[25323]= -720088517;
assign addr[25324]= -791679244;
assign addr[25325]= -862265664;
assign addr[25326]= -931758235;
assign addr[25327]= -1000068799;
assign addr[25328]= -1067110699;
assign addr[25329]= -1132798888;
assign addr[25330]= -1197050035;
assign addr[25331]= -1259782632;
assign addr[25332]= -1320917099;
assign addr[25333]= -1380375881;
assign addr[25334]= -1438083551;
assign addr[25335]= -1493966902;
assign addr[25336]= -1547955041;
assign addr[25337]= -1599979481;
assign addr[25338]= -1649974225;
assign addr[25339]= -1697875851;
assign addr[25340]= -1743623590;
assign addr[25341]= -1787159411;
assign addr[25342]= -1828428082;
assign addr[25343]= -1867377253;
assign addr[25344]= -1903957513;
assign addr[25345]= -1938122457;
assign addr[25346]= -1969828744;
assign addr[25347]= -1999036154;
assign addr[25348]= -2025707632;
assign addr[25349]= -2049809346;
assign addr[25350]= -2071310720;
assign addr[25351]= -2090184478;
assign addr[25352]= -2106406677;
assign addr[25353]= -2119956737;
assign addr[25354]= -2130817471;
assign addr[25355]= -2138975100;
assign addr[25356]= -2144419275;
assign addr[25357]= -2147143090;
assign addr[25358]= -2147143090;
assign addr[25359]= -2144419275;
assign addr[25360]= -2138975100;
assign addr[25361]= -2130817471;
assign addr[25362]= -2119956737;
assign addr[25363]= -2106406677;
assign addr[25364]= -2090184478;
assign addr[25365]= -2071310720;
assign addr[25366]= -2049809346;
assign addr[25367]= -2025707632;
assign addr[25368]= -1999036154;
assign addr[25369]= -1969828744;
assign addr[25370]= -1938122457;
assign addr[25371]= -1903957513;
assign addr[25372]= -1867377253;
assign addr[25373]= -1828428082;
assign addr[25374]= -1787159411;
assign addr[25375]= -1743623590;
assign addr[25376]= -1697875851;
assign addr[25377]= -1649974225;
assign addr[25378]= -1599979481;
assign addr[25379]= -1547955041;
assign addr[25380]= -1493966902;
assign addr[25381]= -1438083551;
assign addr[25382]= -1380375881;
assign addr[25383]= -1320917099;
assign addr[25384]= -1259782632;
assign addr[25385]= -1197050035;
assign addr[25386]= -1132798888;
assign addr[25387]= -1067110699;
assign addr[25388]= -1000068799;
assign addr[25389]= -931758235;
assign addr[25390]= -862265664;
assign addr[25391]= -791679244;
assign addr[25392]= -720088517;
assign addr[25393]= -647584304;
assign addr[25394]= -574258580;
assign addr[25395]= -500204365;
assign addr[25396]= -425515602;
assign addr[25397]= -350287041;
assign addr[25398]= -274614114;
assign addr[25399]= -198592817;
assign addr[25400]= -122319591;
assign addr[25401]= -45891193;
assign addr[25402]= 30595422;
assign addr[25403]= 107043224;
assign addr[25404]= 183355234;
assign addr[25405]= 259434643;
assign addr[25406]= 335184940;
assign addr[25407]= 410510029;
assign addr[25408]= 485314355;
assign addr[25409]= 559503022;
assign addr[25410]= 632981917;
assign addr[25411]= 705657826;
assign addr[25412]= 777438554;
assign addr[25413]= 848233042;
assign addr[25414]= 917951481;
assign addr[25415]= 986505429;
assign addr[25416]= 1053807919;
assign addr[25417]= 1119773573;
assign addr[25418]= 1184318708;
assign addr[25419]= 1247361445;
assign addr[25420]= 1308821808;
assign addr[25421]= 1368621831;
assign addr[25422]= 1426685652;
assign addr[25423]= 1482939614;
assign addr[25424]= 1537312353;
assign addr[25425]= 1589734894;
assign addr[25426]= 1640140734;
assign addr[25427]= 1688465931;
assign addr[25428]= 1734649179;
assign addr[25429]= 1778631892;
assign addr[25430]= 1820358275;
assign addr[25431]= 1859775393;
assign addr[25432]= 1896833245;
assign addr[25433]= 1931484818;
assign addr[25434]= 1963686155;
assign addr[25435]= 1993396407;
assign addr[25436]= 2020577882;
assign addr[25437]= 2045196100;
assign addr[25438]= 2067219829;
assign addr[25439]= 2086621133;
assign addr[25440]= 2103375398;
assign addr[25441]= 2117461370;
assign addr[25442]= 2128861181;
assign addr[25443]= 2137560369;
assign addr[25444]= 2143547897;
assign addr[25445]= 2146816171;
assign addr[25446]= 2147361045;
assign addr[25447]= 2145181827;
assign addr[25448]= 2140281282;
assign addr[25449]= 2132665626;
assign addr[25450]= 2122344521;
assign addr[25451]= 2109331059;
assign addr[25452]= 2093641749;
assign addr[25453]= 2075296495;
assign addr[25454]= 2054318569;
assign addr[25455]= 2030734582;
assign addr[25456]= 2004574453;
assign addr[25457]= 1975871368;
assign addr[25458]= 1944661739;
assign addr[25459]= 1910985158;
assign addr[25460]= 1874884346;
assign addr[25461]= 1836405100;
assign addr[25462]= 1795596234;
assign addr[25463]= 1752509516;
assign addr[25464]= 1707199606;
assign addr[25465]= 1659723983;
assign addr[25466]= 1610142873;
assign addr[25467]= 1558519173;
assign addr[25468]= 1504918373;
assign addr[25469]= 1449408469;
assign addr[25470]= 1392059879;
assign addr[25471]= 1332945355;
assign addr[25472]= 1272139887;
assign addr[25473]= 1209720613;
assign addr[25474]= 1145766716;
assign addr[25475]= 1080359326;
assign addr[25476]= 1013581418;
assign addr[25477]= 945517704;
assign addr[25478]= 876254528;
assign addr[25479]= 805879757;
assign addr[25480]= 734482665;
assign addr[25481]= 662153826;
assign addr[25482]= 588984994;
assign addr[25483]= 515068990;
assign addr[25484]= 440499581;
assign addr[25485]= 365371365;
assign addr[25486]= 289779648;
assign addr[25487]= 213820322;
assign addr[25488]= 137589750;
assign addr[25489]= 61184634;
assign addr[25490]= -15298099;
assign addr[25491]= -91761426;
assign addr[25492]= -168108346;
assign addr[25493]= -244242007;
assign addr[25494]= -320065829;
assign addr[25495]= -395483624;
assign addr[25496]= -470399716;
assign addr[25497]= -544719071;
assign addr[25498]= -618347408;
assign addr[25499]= -691191324;
assign addr[25500]= -763158411;
assign addr[25501]= -834157373;
assign addr[25502]= -904098143;
assign addr[25503]= -972891995;
assign addr[25504]= -1040451659;
assign addr[25505]= -1106691431;
assign addr[25506]= -1171527280;
assign addr[25507]= -1234876957;
assign addr[25508]= -1296660098;
assign addr[25509]= -1356798326;
assign addr[25510]= -1415215352;
assign addr[25511]= -1471837070;
assign addr[25512]= -1526591649;
assign addr[25513]= -1579409630;
assign addr[25514]= -1630224009;
assign addr[25515]= -1678970324;
assign addr[25516]= -1725586737;
assign addr[25517]= -1770014111;
assign addr[25518]= -1812196087;
assign addr[25519]= -1852079154;
assign addr[25520]= -1889612716;
assign addr[25521]= -1924749160;
assign addr[25522]= -1957443913;
assign addr[25523]= -1987655498;
assign addr[25524]= -2015345591;
assign addr[25525]= -2040479063;
assign addr[25526]= -2063024031;
assign addr[25527]= -2082951896;
assign addr[25528]= -2100237377;
assign addr[25529]= -2114858546;
assign addr[25530]= -2126796855;
assign addr[25531]= -2136037160;
assign addr[25532]= -2142567738;
assign addr[25533]= -2146380306;
assign addr[25534]= -2147470025;
assign addr[25535]= -2145835515;
assign addr[25536]= -2141478848;
assign addr[25537]= -2134405552;
assign addr[25538]= -2124624598;
assign addr[25539]= -2112148396;
assign addr[25540]= -2096992772;
assign addr[25541]= -2079176953;
assign addr[25542]= -2058723538;
assign addr[25543]= -2035658475;
assign addr[25544]= -2010011024;
assign addr[25545]= -1981813720;
assign addr[25546]= -1951102334;
assign addr[25547]= -1917915825;
assign addr[25548]= -1882296293;
assign addr[25549]= -1844288924;
assign addr[25550]= -1803941934;
assign addr[25551]= -1761306505;
assign addr[25552]= -1716436725;
assign addr[25553]= -1669389513;
assign addr[25554]= -1620224553;
assign addr[25555]= -1569004214;
assign addr[25556]= -1515793473;
assign addr[25557]= -1460659832;
assign addr[25558]= -1403673233;
assign addr[25559]= -1344905966;
assign addr[25560]= -1284432584;
assign addr[25561]= -1222329801;
assign addr[25562]= -1158676398;
assign addr[25563]= -1093553126;
assign addr[25564]= -1027042599;
assign addr[25565]= -959229189;
assign addr[25566]= -890198924;
assign addr[25567]= -820039373;
assign addr[25568]= -748839539;
assign addr[25569]= -676689746;
assign addr[25570]= -603681519;
assign addr[25571]= -529907477;
assign addr[25572]= -455461206;
assign addr[25573]= -380437148;
assign addr[25574]= -304930476;
assign addr[25575]= -229036977;
assign addr[25576]= -152852926;
assign addr[25577]= -76474970;
assign addr[25578]= 0;
assign addr[25579]= 76474970;
assign addr[25580]= 152852926;
assign addr[25581]= 229036977;
assign addr[25582]= 304930476;
assign addr[25583]= 380437148;
assign addr[25584]= 455461206;
assign addr[25585]= 529907477;
assign addr[25586]= 603681519;
assign addr[25587]= 676689746;
assign addr[25588]= 748839539;
assign addr[25589]= 820039373;
assign addr[25590]= 890198924;
assign addr[25591]= 959229189;
assign addr[25592]= 1027042599;
assign addr[25593]= 1093553126;
assign addr[25594]= 1158676398;
assign addr[25595]= 1222329801;
assign addr[25596]= 1284432584;
assign addr[25597]= 1344905966;
assign addr[25598]= 1403673233;
assign addr[25599]= 1460659832;
assign addr[25600]= 1515793473;
assign addr[25601]= 1569004214;
assign addr[25602]= 1620224553;
assign addr[25603]= 1669389513;
assign addr[25604]= 1716436725;
assign addr[25605]= 1761306505;
assign addr[25606]= 1803941934;
assign addr[25607]= 1844288924;
assign addr[25608]= 1882296293;
assign addr[25609]= 1917915825;
assign addr[25610]= 1951102334;
assign addr[25611]= 1981813720;
assign addr[25612]= 2010011024;
assign addr[25613]= 2035658475;
assign addr[25614]= 2058723538;
assign addr[25615]= 2079176953;
assign addr[25616]= 2096992772;
assign addr[25617]= 2112148396;
assign addr[25618]= 2124624598;
assign addr[25619]= 2134405552;
assign addr[25620]= 2141478848;
assign addr[25621]= 2145835515;
assign addr[25622]= 2147470025;
assign addr[25623]= 2146380306;
assign addr[25624]= 2142567738;
assign addr[25625]= 2136037160;
assign addr[25626]= 2126796855;
assign addr[25627]= 2114858546;
assign addr[25628]= 2100237377;
assign addr[25629]= 2082951896;
assign addr[25630]= 2063024031;
assign addr[25631]= 2040479063;
assign addr[25632]= 2015345591;
assign addr[25633]= 1987655498;
assign addr[25634]= 1957443913;
assign addr[25635]= 1924749160;
assign addr[25636]= 1889612716;
assign addr[25637]= 1852079154;
assign addr[25638]= 1812196087;
assign addr[25639]= 1770014111;
assign addr[25640]= 1725586737;
assign addr[25641]= 1678970324;
assign addr[25642]= 1630224009;
assign addr[25643]= 1579409630;
assign addr[25644]= 1526591649;
assign addr[25645]= 1471837070;
assign addr[25646]= 1415215352;
assign addr[25647]= 1356798326;
assign addr[25648]= 1296660098;
assign addr[25649]= 1234876957;
assign addr[25650]= 1171527280;
assign addr[25651]= 1106691431;
assign addr[25652]= 1040451659;
assign addr[25653]= 972891995;
assign addr[25654]= 904098143;
assign addr[25655]= 834157373;
assign addr[25656]= 763158411;
assign addr[25657]= 691191324;
assign addr[25658]= 618347408;
assign addr[25659]= 544719071;
assign addr[25660]= 470399716;
assign addr[25661]= 395483624;
assign addr[25662]= 320065829;
assign addr[25663]= 244242007;
assign addr[25664]= 168108346;
assign addr[25665]= 91761426;
assign addr[25666]= 15298099;
assign addr[25667]= -61184634;
assign addr[25668]= -137589750;
assign addr[25669]= -213820322;
assign addr[25670]= -289779648;
assign addr[25671]= -365371365;
assign addr[25672]= -440499581;
assign addr[25673]= -515068990;
assign addr[25674]= -588984994;
assign addr[25675]= -662153826;
assign addr[25676]= -734482665;
assign addr[25677]= -805879757;
assign addr[25678]= -876254528;
assign addr[25679]= -945517704;
assign addr[25680]= -1013581418;
assign addr[25681]= -1080359326;
assign addr[25682]= -1145766716;
assign addr[25683]= -1209720613;
assign addr[25684]= -1272139887;
assign addr[25685]= -1332945355;
assign addr[25686]= -1392059879;
assign addr[25687]= -1449408469;
assign addr[25688]= -1504918373;
assign addr[25689]= -1558519173;
assign addr[25690]= -1610142873;
assign addr[25691]= -1659723983;
assign addr[25692]= -1707199606;
assign addr[25693]= -1752509516;
assign addr[25694]= -1795596234;
assign addr[25695]= -1836405100;
assign addr[25696]= -1874884346;
assign addr[25697]= -1910985158;
assign addr[25698]= -1944661739;
assign addr[25699]= -1975871368;
assign addr[25700]= -2004574453;
assign addr[25701]= -2030734582;
assign addr[25702]= -2054318569;
assign addr[25703]= -2075296495;
assign addr[25704]= -2093641749;
assign addr[25705]= -2109331059;
assign addr[25706]= -2122344521;
assign addr[25707]= -2132665626;
assign addr[25708]= -2140281282;
assign addr[25709]= -2145181827;
assign addr[25710]= -2147361045;
assign addr[25711]= -2146816171;
assign addr[25712]= -2143547897;
assign addr[25713]= -2137560369;
assign addr[25714]= -2128861181;
assign addr[25715]= -2117461370;
assign addr[25716]= -2103375398;
assign addr[25717]= -2086621133;
assign addr[25718]= -2067219829;
assign addr[25719]= -2045196100;
assign addr[25720]= -2020577882;
assign addr[25721]= -1993396407;
assign addr[25722]= -1963686155;
assign addr[25723]= -1931484818;
assign addr[25724]= -1896833245;
assign addr[25725]= -1859775393;
assign addr[25726]= -1820358275;
assign addr[25727]= -1778631892;
assign addr[25728]= -1734649179;
assign addr[25729]= -1688465931;
assign addr[25730]= -1640140734;
assign addr[25731]= -1589734894;
assign addr[25732]= -1537312353;
assign addr[25733]= -1482939614;
assign addr[25734]= -1426685652;
assign addr[25735]= -1368621831;
assign addr[25736]= -1308821808;
assign addr[25737]= -1247361445;
assign addr[25738]= -1184318708;
assign addr[25739]= -1119773573;
assign addr[25740]= -1053807919;
assign addr[25741]= -986505429;
assign addr[25742]= -917951481;
assign addr[25743]= -848233042;
assign addr[25744]= -777438554;
assign addr[25745]= -705657826;
assign addr[25746]= -632981917;
assign addr[25747]= -559503022;
assign addr[25748]= -485314355;
assign addr[25749]= -410510029;
assign addr[25750]= -335184940;
assign addr[25751]= -259434643;
assign addr[25752]= -183355234;
assign addr[25753]= -107043224;
assign addr[25754]= -30595422;
assign addr[25755]= 45891193;
assign addr[25756]= 122319591;
assign addr[25757]= 198592817;
assign addr[25758]= 274614114;
assign addr[25759]= 350287041;
assign addr[25760]= 425515602;
assign addr[25761]= 500204365;
assign addr[25762]= 574258580;
assign addr[25763]= 647584304;
assign addr[25764]= 720088517;
assign addr[25765]= 791679244;
assign addr[25766]= 862265664;
assign addr[25767]= 931758235;
assign addr[25768]= 1000068799;
assign addr[25769]= 1067110699;
assign addr[25770]= 1132798888;
assign addr[25771]= 1197050035;
assign addr[25772]= 1259782632;
assign addr[25773]= 1320917099;
assign addr[25774]= 1380375881;
assign addr[25775]= 1438083551;
assign addr[25776]= 1493966902;
assign addr[25777]= 1547955041;
assign addr[25778]= 1599979481;
assign addr[25779]= 1649974225;
assign addr[25780]= 1697875851;
assign addr[25781]= 1743623590;
assign addr[25782]= 1787159411;
assign addr[25783]= 1828428082;
assign addr[25784]= 1867377253;
assign addr[25785]= 1903957513;
assign addr[25786]= 1938122457;
assign addr[25787]= 1969828744;
assign addr[25788]= 1999036154;
assign addr[25789]= 2025707632;
assign addr[25790]= 2049809346;
assign addr[25791]= 2071310720;
assign addr[25792]= 2090184478;
assign addr[25793]= 2106406677;
assign addr[25794]= 2119956737;
assign addr[25795]= 2130817471;
assign addr[25796]= 2138975100;
assign addr[25797]= 2144419275;
assign addr[25798]= 2147143090;
assign addr[25799]= 2147143090;
assign addr[25800]= 2144419275;
assign addr[25801]= 2138975100;
assign addr[25802]= 2130817471;
assign addr[25803]= 2119956737;
assign addr[25804]= 2106406677;
assign addr[25805]= 2090184478;
assign addr[25806]= 2071310720;
assign addr[25807]= 2049809346;
assign addr[25808]= 2025707632;
assign addr[25809]= 1999036154;
assign addr[25810]= 1969828744;
assign addr[25811]= 1938122457;
assign addr[25812]= 1903957513;
assign addr[25813]= 1867377253;
assign addr[25814]= 1828428082;
assign addr[25815]= 1787159411;
assign addr[25816]= 1743623590;
assign addr[25817]= 1697875851;
assign addr[25818]= 1649974225;
assign addr[25819]= 1599979481;
assign addr[25820]= 1547955041;
assign addr[25821]= 1493966902;
assign addr[25822]= 1438083551;
assign addr[25823]= 1380375881;
assign addr[25824]= 1320917099;
assign addr[25825]= 1259782632;
assign addr[25826]= 1197050035;
assign addr[25827]= 1132798888;
assign addr[25828]= 1067110699;
assign addr[25829]= 1000068799;
assign addr[25830]= 931758235;
assign addr[25831]= 862265664;
assign addr[25832]= 791679244;
assign addr[25833]= 720088517;
assign addr[25834]= 647584304;
assign addr[25835]= 574258580;
assign addr[25836]= 500204365;
assign addr[25837]= 425515602;
assign addr[25838]= 350287041;
assign addr[25839]= 274614114;
assign addr[25840]= 198592817;
assign addr[25841]= 122319591;
assign addr[25842]= 45891193;
assign addr[25843]= -30595422;
assign addr[25844]= -107043224;
assign addr[25845]= -183355234;
assign addr[25846]= -259434643;
assign addr[25847]= -335184940;
assign addr[25848]= -410510029;
assign addr[25849]= -485314355;
assign addr[25850]= -559503022;
assign addr[25851]= -632981917;
assign addr[25852]= -705657826;
assign addr[25853]= -777438554;
assign addr[25854]= -848233042;
assign addr[25855]= -917951481;
assign addr[25856]= -986505429;
assign addr[25857]= -1053807919;
assign addr[25858]= -1119773573;
assign addr[25859]= -1184318708;
assign addr[25860]= -1247361445;
assign addr[25861]= -1308821808;
assign addr[25862]= -1368621831;
assign addr[25863]= -1426685652;
assign addr[25864]= -1482939614;
assign addr[25865]= -1537312353;
assign addr[25866]= -1589734894;
assign addr[25867]= -1640140734;
assign addr[25868]= -1688465931;
assign addr[25869]= -1734649179;
assign addr[25870]= -1778631892;
assign addr[25871]= -1820358275;
assign addr[25872]= -1859775393;
assign addr[25873]= -1896833245;
assign addr[25874]= -1931484818;
assign addr[25875]= -1963686155;
assign addr[25876]= -1993396407;
assign addr[25877]= -2020577882;
assign addr[25878]= -2045196100;
assign addr[25879]= -2067219829;
assign addr[25880]= -2086621133;
assign addr[25881]= -2103375398;
assign addr[25882]= -2117461370;
assign addr[25883]= -2128861181;
assign addr[25884]= -2137560369;
assign addr[25885]= -2143547897;
assign addr[25886]= -2146816171;
assign addr[25887]= -2147361045;
assign addr[25888]= -2145181827;
assign addr[25889]= -2140281282;
assign addr[25890]= -2132665626;
assign addr[25891]= -2122344521;
assign addr[25892]= -2109331059;
assign addr[25893]= -2093641749;
assign addr[25894]= -2075296495;
assign addr[25895]= -2054318569;
assign addr[25896]= -2030734582;
assign addr[25897]= -2004574453;
assign addr[25898]= -1975871368;
assign addr[25899]= -1944661739;
assign addr[25900]= -1910985158;
assign addr[25901]= -1874884346;
assign addr[25902]= -1836405100;
assign addr[25903]= -1795596234;
assign addr[25904]= -1752509516;
assign addr[25905]= -1707199606;
assign addr[25906]= -1659723983;
assign addr[25907]= -1610142873;
assign addr[25908]= -1558519173;
assign addr[25909]= -1504918373;
assign addr[25910]= -1449408469;
assign addr[25911]= -1392059879;
assign addr[25912]= -1332945355;
assign addr[25913]= -1272139887;
assign addr[25914]= -1209720613;
assign addr[25915]= -1145766716;
assign addr[25916]= -1080359326;
assign addr[25917]= -1013581418;
assign addr[25918]= -945517704;
assign addr[25919]= -876254528;
assign addr[25920]= -805879757;
assign addr[25921]= -734482665;
assign addr[25922]= -662153826;
assign addr[25923]= -588984994;
assign addr[25924]= -515068990;
assign addr[25925]= -440499581;
assign addr[25926]= -365371365;
assign addr[25927]= -289779648;
assign addr[25928]= -213820322;
assign addr[25929]= -137589750;
assign addr[25930]= -61184634;
assign addr[25931]= 15298099;
assign addr[25932]= 91761426;
assign addr[25933]= 168108346;
assign addr[25934]= 244242007;
assign addr[25935]= 320065829;
assign addr[25936]= 395483624;
assign addr[25937]= 470399716;
assign addr[25938]= 544719071;
assign addr[25939]= 618347408;
assign addr[25940]= 691191324;
assign addr[25941]= 763158411;
assign addr[25942]= 834157373;
assign addr[25943]= 904098143;
assign addr[25944]= 972891995;
assign addr[25945]= 1040451659;
assign addr[25946]= 1106691431;
assign addr[25947]= 1171527280;
assign addr[25948]= 1234876957;
assign addr[25949]= 1296660098;
assign addr[25950]= 1356798326;
assign addr[25951]= 1415215352;
assign addr[25952]= 1471837070;
assign addr[25953]= 1526591649;
assign addr[25954]= 1579409630;
assign addr[25955]= 1630224009;
assign addr[25956]= 1678970324;
assign addr[25957]= 1725586737;
assign addr[25958]= 1770014111;
assign addr[25959]= 1812196087;
assign addr[25960]= 1852079154;
assign addr[25961]= 1889612716;
assign addr[25962]= 1924749160;
assign addr[25963]= 1957443913;
assign addr[25964]= 1987655498;
assign addr[25965]= 2015345591;
assign addr[25966]= 2040479063;
assign addr[25967]= 2063024031;
assign addr[25968]= 2082951896;
assign addr[25969]= 2100237377;
assign addr[25970]= 2114858546;
assign addr[25971]= 2126796855;
assign addr[25972]= 2136037160;
assign addr[25973]= 2142567738;
assign addr[25974]= 2146380306;
assign addr[25975]= 2147470025;
assign addr[25976]= 2145835515;
assign addr[25977]= 2141478848;
assign addr[25978]= 2134405552;
assign addr[25979]= 2124624598;
assign addr[25980]= 2112148396;
assign addr[25981]= 2096992772;
assign addr[25982]= 2079176953;
assign addr[25983]= 2058723538;
assign addr[25984]= 2035658475;
assign addr[25985]= 2010011024;
assign addr[25986]= 1981813720;
assign addr[25987]= 1951102334;
assign addr[25988]= 1917915825;
assign addr[25989]= 1882296293;
assign addr[25990]= 1844288924;
assign addr[25991]= 1803941934;
assign addr[25992]= 1761306505;
assign addr[25993]= 1716436725;
assign addr[25994]= 1669389513;
assign addr[25995]= 1620224553;
assign addr[25996]= 1569004214;
assign addr[25997]= 1515793473;
assign addr[25998]= 1460659832;
assign addr[25999]= 1403673233;
assign addr[26000]= 1344905966;
assign addr[26001]= 1284432584;
assign addr[26002]= 1222329801;
assign addr[26003]= 1158676398;
assign addr[26004]= 1093553126;
assign addr[26005]= 1027042599;
assign addr[26006]= 959229189;
assign addr[26007]= 890198924;
assign addr[26008]= 820039373;
assign addr[26009]= 748839539;
assign addr[26010]= 676689746;
assign addr[26011]= 603681519;
assign addr[26012]= 529907477;
assign addr[26013]= 455461206;
assign addr[26014]= 380437148;
assign addr[26015]= 304930476;
assign addr[26016]= 229036977;
assign addr[26017]= 152852926;
assign addr[26018]= 76474970;
assign addr[26019]= 0;
assign addr[26020]= -76474970;
assign addr[26021]= -152852926;
assign addr[26022]= -229036977;
assign addr[26023]= -304930476;
assign addr[26024]= -380437148;
assign addr[26025]= -455461206;
assign addr[26026]= -529907477;
assign addr[26027]= -603681519;
assign addr[26028]= -676689746;
assign addr[26029]= -748839539;
assign addr[26030]= -820039373;
assign addr[26031]= -890198924;
assign addr[26032]= -959229189;
assign addr[26033]= -1027042599;
assign addr[26034]= -1093553126;
assign addr[26035]= -1158676398;
assign addr[26036]= -1222329801;
assign addr[26037]= -1284432584;
assign addr[26038]= -1344905966;
assign addr[26039]= -1403673233;
assign addr[26040]= -1460659832;
assign addr[26041]= -1515793473;
assign addr[26042]= -1569004214;
assign addr[26043]= -1620224553;
assign addr[26044]= -1669389513;
assign addr[26045]= -1716436725;
assign addr[26046]= -1761306505;
assign addr[26047]= -1803941934;
assign addr[26048]= -1844288924;
assign addr[26049]= -1882296293;
assign addr[26050]= -1917915825;
assign addr[26051]= -1951102334;
assign addr[26052]= -1981813720;
assign addr[26053]= -2010011024;
assign addr[26054]= -2035658475;
assign addr[26055]= -2058723538;
assign addr[26056]= -2079176953;
assign addr[26057]= -2096992772;
assign addr[26058]= -2112148396;
assign addr[26059]= -2124624598;
assign addr[26060]= -2134405552;
assign addr[26061]= -2141478848;
assign addr[26062]= -2145835515;
assign addr[26063]= -2147470025;
assign addr[26064]= -2146380306;
assign addr[26065]= -2142567738;
assign addr[26066]= -2136037160;
assign addr[26067]= -2126796855;
assign addr[26068]= -2114858546;
assign addr[26069]= -2100237377;
assign addr[26070]= -2082951896;
assign addr[26071]= -2063024031;
assign addr[26072]= -2040479063;
assign addr[26073]= -2015345591;
assign addr[26074]= -1987655498;
assign addr[26075]= -1957443913;
assign addr[26076]= -1924749160;
assign addr[26077]= -1889612716;
assign addr[26078]= -1852079154;
assign addr[26079]= -1812196087;
assign addr[26080]= -1770014111;
assign addr[26081]= -1725586737;
assign addr[26082]= -1678970324;
assign addr[26083]= -1630224009;
assign addr[26084]= -1579409630;
assign addr[26085]= -1526591649;
assign addr[26086]= -1471837070;
assign addr[26087]= -1415215352;
assign addr[26088]= -1356798326;
assign addr[26089]= -1296660098;
assign addr[26090]= -1234876957;
assign addr[26091]= -1171527280;
assign addr[26092]= -1106691431;
assign addr[26093]= -1040451659;
assign addr[26094]= -972891995;
assign addr[26095]= -904098143;
assign addr[26096]= -834157373;
assign addr[26097]= -763158411;
assign addr[26098]= -691191324;
assign addr[26099]= -618347408;
assign addr[26100]= -544719071;
assign addr[26101]= -470399716;
assign addr[26102]= -395483624;
assign addr[26103]= -320065829;
assign addr[26104]= -244242007;
assign addr[26105]= -168108346;
assign addr[26106]= -91761426;
assign addr[26107]= -15298099;
assign addr[26108]= 61184634;
assign addr[26109]= 137589750;
assign addr[26110]= 213820322;
assign addr[26111]= 289779648;
assign addr[26112]= 365371365;
assign addr[26113]= 440499581;
assign addr[26114]= 515068990;
assign addr[26115]= 588984994;
assign addr[26116]= 662153826;
assign addr[26117]= 734482665;
assign addr[26118]= 805879757;
assign addr[26119]= 876254528;
assign addr[26120]= 945517704;
assign addr[26121]= 1013581418;
assign addr[26122]= 1080359326;
assign addr[26123]= 1145766716;
assign addr[26124]= 1209720613;
assign addr[26125]= 1272139887;
assign addr[26126]= 1332945355;
assign addr[26127]= 1392059879;
assign addr[26128]= 1449408469;
assign addr[26129]= 1504918373;
assign addr[26130]= 1558519173;
assign addr[26131]= 1610142873;
assign addr[26132]= 1659723983;
assign addr[26133]= 1707199606;
assign addr[26134]= 1752509516;
assign addr[26135]= 1795596234;
assign addr[26136]= 1836405100;
assign addr[26137]= 1874884346;
assign addr[26138]= 1910985158;
assign addr[26139]= 1944661739;
assign addr[26140]= 1975871368;
assign addr[26141]= 2004574453;
assign addr[26142]= 2030734582;
assign addr[26143]= 2054318569;
assign addr[26144]= 2075296495;
assign addr[26145]= 2093641749;
assign addr[26146]= 2109331059;
assign addr[26147]= 2122344521;
assign addr[26148]= 2132665626;
assign addr[26149]= 2140281282;
assign addr[26150]= 2145181827;
assign addr[26151]= 2147361045;
assign addr[26152]= 2146816171;
assign addr[26153]= 2143547897;
assign addr[26154]= 2137560369;
assign addr[26155]= 2128861181;
assign addr[26156]= 2117461370;
assign addr[26157]= 2103375398;
assign addr[26158]= 2086621133;
assign addr[26159]= 2067219829;
assign addr[26160]= 2045196100;
assign addr[26161]= 2020577882;
assign addr[26162]= 1993396407;
assign addr[26163]= 1963686155;
assign addr[26164]= 1931484818;
assign addr[26165]= 1896833245;
assign addr[26166]= 1859775393;
assign addr[26167]= 1820358275;
assign addr[26168]= 1778631892;
assign addr[26169]= 1734649179;
assign addr[26170]= 1688465931;
assign addr[26171]= 1640140734;
assign addr[26172]= 1589734894;
assign addr[26173]= 1537312353;
assign addr[26174]= 1482939614;
assign addr[26175]= 1426685652;
assign addr[26176]= 1368621831;
assign addr[26177]= 1308821808;
assign addr[26178]= 1247361445;
assign addr[26179]= 1184318708;
assign addr[26180]= 1119773573;
assign addr[26181]= 1053807919;
assign addr[26182]= 986505429;
assign addr[26183]= 917951481;
assign addr[26184]= 848233042;
assign addr[26185]= 777438554;
assign addr[26186]= 705657826;
assign addr[26187]= 632981917;
assign addr[26188]= 559503022;
assign addr[26189]= 485314355;
assign addr[26190]= 410510029;
assign addr[26191]= 335184940;
assign addr[26192]= 259434643;
assign addr[26193]= 183355234;
assign addr[26194]= 107043224;
assign addr[26195]= 30595422;
assign addr[26196]= -45891193;
assign addr[26197]= -122319591;
assign addr[26198]= -198592817;
assign addr[26199]= -274614114;
assign addr[26200]= -350287041;
assign addr[26201]= -425515602;
assign addr[26202]= -500204365;
assign addr[26203]= -574258580;
assign addr[26204]= -647584304;
assign addr[26205]= -720088517;
assign addr[26206]= -791679244;
assign addr[26207]= -862265664;
assign addr[26208]= -931758235;
assign addr[26209]= -1000068799;
assign addr[26210]= -1067110699;
assign addr[26211]= -1132798888;
assign addr[26212]= -1197050035;
assign addr[26213]= -1259782632;
assign addr[26214]= -1320917099;
assign addr[26215]= -1380375881;
assign addr[26216]= -1438083551;
assign addr[26217]= -1493966902;
assign addr[26218]= -1547955041;
assign addr[26219]= -1599979481;
assign addr[26220]= -1649974225;
assign addr[26221]= -1697875851;
assign addr[26222]= -1743623590;
assign addr[26223]= -1787159411;
assign addr[26224]= -1828428082;
assign addr[26225]= -1867377253;
assign addr[26226]= -1903957513;
assign addr[26227]= -1938122457;
assign addr[26228]= -1969828744;
assign addr[26229]= -1999036154;
assign addr[26230]= -2025707632;
assign addr[26231]= -2049809346;
assign addr[26232]= -2071310720;
assign addr[26233]= -2090184478;
assign addr[26234]= -2106406677;
assign addr[26235]= -2119956737;
assign addr[26236]= -2130817471;
assign addr[26237]= -2138975100;
assign addr[26238]= -2144419275;
assign addr[26239]= -2147143090;
assign addr[26240]= -2147143090;
assign addr[26241]= -2144419275;
assign addr[26242]= -2138975100;
assign addr[26243]= -2130817471;
assign addr[26244]= -2119956737;
assign addr[26245]= -2106406677;
assign addr[26246]= -2090184478;
assign addr[26247]= -2071310720;
assign addr[26248]= -2049809346;
assign addr[26249]= -2025707632;
assign addr[26250]= -1999036154;
assign addr[26251]= -1969828744;
assign addr[26252]= -1938122457;
assign addr[26253]= -1903957513;
assign addr[26254]= -1867377253;
assign addr[26255]= -1828428082;
assign addr[26256]= -1787159411;
assign addr[26257]= -1743623590;
assign addr[26258]= -1697875851;
assign addr[26259]= -1649974225;
assign addr[26260]= -1599979481;
assign addr[26261]= -1547955041;
assign addr[26262]= -1493966902;
assign addr[26263]= -1438083551;
assign addr[26264]= -1380375881;
assign addr[26265]= -1320917099;
assign addr[26266]= -1259782632;
assign addr[26267]= -1197050035;
assign addr[26268]= -1132798888;
assign addr[26269]= -1067110699;
assign addr[26270]= -1000068799;
assign addr[26271]= -931758235;
assign addr[26272]= -862265664;
assign addr[26273]= -791679244;
assign addr[26274]= -720088517;
assign addr[26275]= -647584304;
assign addr[26276]= -574258580;
assign addr[26277]= -500204365;
assign addr[26278]= -425515602;
assign addr[26279]= -350287041;
assign addr[26280]= -274614114;
assign addr[26281]= -198592817;
assign addr[26282]= -122319591;
assign addr[26283]= -45891193;
assign addr[26284]= 30595422;
assign addr[26285]= 107043224;
assign addr[26286]= 183355234;
assign addr[26287]= 259434643;
assign addr[26288]= 335184940;
assign addr[26289]= 410510029;
assign addr[26290]= 485314355;
assign addr[26291]= 559503022;
assign addr[26292]= 632981917;
assign addr[26293]= 705657826;
assign addr[26294]= 777438554;
assign addr[26295]= 848233042;
assign addr[26296]= 917951481;
assign addr[26297]= 986505429;
assign addr[26298]= 1053807919;
assign addr[26299]= 1119773573;
assign addr[26300]= 1184318708;
assign addr[26301]= 1247361445;
assign addr[26302]= 1308821808;
assign addr[26303]= 1368621831;
assign addr[26304]= 1426685652;
assign addr[26305]= 1482939614;
assign addr[26306]= 1537312353;
assign addr[26307]= 1589734894;
assign addr[26308]= 1640140734;
assign addr[26309]= 1688465931;
assign addr[26310]= 1734649179;
assign addr[26311]= 1778631892;
assign addr[26312]= 1820358275;
assign addr[26313]= 1859775393;
assign addr[26314]= 1896833245;
assign addr[26315]= 1931484818;
assign addr[26316]= 1963686155;
assign addr[26317]= 1993396407;
assign addr[26318]= 2020577882;
assign addr[26319]= 2045196100;
assign addr[26320]= 2067219829;
assign addr[26321]= 2086621133;
assign addr[26322]= 2103375398;
assign addr[26323]= 2117461370;
assign addr[26324]= 2128861181;
assign addr[26325]= 2137560369;
assign addr[26326]= 2143547897;
assign addr[26327]= 2146816171;
assign addr[26328]= 2147361045;
assign addr[26329]= 2145181827;
assign addr[26330]= 2140281282;
assign addr[26331]= 2132665626;
assign addr[26332]= 2122344521;
assign addr[26333]= 2109331059;
assign addr[26334]= 2093641749;
assign addr[26335]= 2075296495;
assign addr[26336]= 2054318569;
assign addr[26337]= 2030734582;
assign addr[26338]= 2004574453;
assign addr[26339]= 1975871368;
assign addr[26340]= 1944661739;
assign addr[26341]= 1910985158;
assign addr[26342]= 1874884346;
assign addr[26343]= 1836405100;
assign addr[26344]= 1795596234;
assign addr[26345]= 1752509516;
assign addr[26346]= 1707199606;
assign addr[26347]= 1659723983;
assign addr[26348]= 1610142873;
assign addr[26349]= 1558519173;
assign addr[26350]= 1504918373;
assign addr[26351]= 1449408469;
assign addr[26352]= 1392059879;
assign addr[26353]= 1332945355;
assign addr[26354]= 1272139887;
assign addr[26355]= 1209720613;
assign addr[26356]= 1145766716;
assign addr[26357]= 1080359326;
assign addr[26358]= 1013581418;
assign addr[26359]= 945517704;
assign addr[26360]= 876254528;
assign addr[26361]= 805879757;
assign addr[26362]= 734482665;
assign addr[26363]= 662153826;
assign addr[26364]= 588984994;
assign addr[26365]= 515068990;
assign addr[26366]= 440499581;
assign addr[26367]= 365371365;
assign addr[26368]= 289779648;
assign addr[26369]= 213820322;
assign addr[26370]= 137589750;
assign addr[26371]= 61184634;
assign addr[26372]= -15298099;
assign addr[26373]= -91761426;
assign addr[26374]= -168108346;
assign addr[26375]= -244242007;
assign addr[26376]= -320065829;
assign addr[26377]= -395483624;
assign addr[26378]= -470399716;
assign addr[26379]= -544719071;
assign addr[26380]= -618347408;
assign addr[26381]= -691191324;
assign addr[26382]= -763158411;
assign addr[26383]= -834157373;
assign addr[26384]= -904098143;
assign addr[26385]= -972891995;
assign addr[26386]= -1040451659;
assign addr[26387]= -1106691431;
assign addr[26388]= -1171527280;
assign addr[26389]= -1234876957;
assign addr[26390]= -1296660098;
assign addr[26391]= -1356798326;
assign addr[26392]= -1415215352;
assign addr[26393]= -1471837070;
assign addr[26394]= -1526591649;
assign addr[26395]= -1579409630;
assign addr[26396]= -1630224009;
assign addr[26397]= -1678970324;
assign addr[26398]= -1725586737;
assign addr[26399]= -1770014111;
assign addr[26400]= -1812196087;
assign addr[26401]= -1852079154;
assign addr[26402]= -1889612716;
assign addr[26403]= -1924749160;
assign addr[26404]= -1957443913;
assign addr[26405]= -1987655498;
assign addr[26406]= -2015345591;
assign addr[26407]= -2040479063;
assign addr[26408]= -2063024031;
assign addr[26409]= -2082951896;
assign addr[26410]= -2100237377;
assign addr[26411]= -2114858546;
assign addr[26412]= -2126796855;
assign addr[26413]= -2136037160;
assign addr[26414]= -2142567738;
assign addr[26415]= -2146380306;
assign addr[26416]= -2147470025;
assign addr[26417]= -2145835515;
assign addr[26418]= -2141478848;
assign addr[26419]= -2134405552;
assign addr[26420]= -2124624598;
assign addr[26421]= -2112148396;
assign addr[26422]= -2096992772;
assign addr[26423]= -2079176953;
assign addr[26424]= -2058723538;
assign addr[26425]= -2035658475;
assign addr[26426]= -2010011024;
assign addr[26427]= -1981813720;
assign addr[26428]= -1951102334;
assign addr[26429]= -1917915825;
assign addr[26430]= -1882296293;
assign addr[26431]= -1844288924;
assign addr[26432]= -1803941934;
assign addr[26433]= -1761306505;
assign addr[26434]= -1716436725;
assign addr[26435]= -1669389513;
assign addr[26436]= -1620224553;
assign addr[26437]= -1569004214;
assign addr[26438]= -1515793473;
assign addr[26439]= -1460659832;
assign addr[26440]= -1403673233;
assign addr[26441]= -1344905966;
assign addr[26442]= -1284432584;
assign addr[26443]= -1222329801;
assign addr[26444]= -1158676398;
assign addr[26445]= -1093553126;
assign addr[26446]= -1027042599;
assign addr[26447]= -959229189;
assign addr[26448]= -890198924;
assign addr[26449]= -820039373;
assign addr[26450]= -748839539;
assign addr[26451]= -676689746;
assign addr[26452]= -603681519;
assign addr[26453]= -529907477;
assign addr[26454]= -455461206;
assign addr[26455]= -380437148;
assign addr[26456]= -304930476;
assign addr[26457]= -229036977;
assign addr[26458]= -152852926;
assign addr[26459]= -76474970;
assign addr[26460]= 0;
assign addr[26461]= 76474970;
assign addr[26462]= 152852926;
assign addr[26463]= 229036977;
assign addr[26464]= 304930476;
assign addr[26465]= 380437148;
assign addr[26466]= 455461206;
assign addr[26467]= 529907477;
assign addr[26468]= 603681519;
assign addr[26469]= 676689746;
assign addr[26470]= 748839539;
assign addr[26471]= 820039373;
assign addr[26472]= 890198924;
assign addr[26473]= 959229189;
assign addr[26474]= 1027042599;
assign addr[26475]= 1093553126;
assign addr[26476]= 1158676398;
assign addr[26477]= 1222329801;
assign addr[26478]= 1284432584;
assign addr[26479]= 1344905966;
assign addr[26480]= 1403673233;
assign addr[26481]= 1460659832;
assign addr[26482]= 1515793473;
assign addr[26483]= 1569004214;
assign addr[26484]= 1620224553;
assign addr[26485]= 1669389513;
assign addr[26486]= 1716436725;
assign addr[26487]= 1761306505;
assign addr[26488]= 1803941934;
assign addr[26489]= 1844288924;
assign addr[26490]= 1882296293;
assign addr[26491]= 1917915825;
assign addr[26492]= 1951102334;
assign addr[26493]= 1981813720;
assign addr[26494]= 2010011024;
assign addr[26495]= 2035658475;
assign addr[26496]= 2058723538;
assign addr[26497]= 2079176953;
assign addr[26498]= 2096992772;
assign addr[26499]= 2112148396;
assign addr[26500]= 2124624598;
assign addr[26501]= 2134405552;
assign addr[26502]= 2141478848;
assign addr[26503]= 2145835515;
assign addr[26504]= 2147470025;
assign addr[26505]= 2146380306;
assign addr[26506]= 2142567738;
assign addr[26507]= 2136037160;
assign addr[26508]= 2126796855;
assign addr[26509]= 2114858546;
assign addr[26510]= 2100237377;
assign addr[26511]= 2082951896;
assign addr[26512]= 2063024031;
assign addr[26513]= 2040479063;
assign addr[26514]= 2015345591;
assign addr[26515]= 1987655498;
assign addr[26516]= 1957443913;
assign addr[26517]= 1924749160;
assign addr[26518]= 1889612716;
assign addr[26519]= 1852079154;
assign addr[26520]= 1812196087;
assign addr[26521]= 1770014111;
assign addr[26522]= 1725586737;
assign addr[26523]= 1678970324;
assign addr[26524]= 1630224009;
assign addr[26525]= 1579409630;
assign addr[26526]= 1526591649;
assign addr[26527]= 1471837070;
assign addr[26528]= 1415215352;
assign addr[26529]= 1356798326;
assign addr[26530]= 1296660098;
assign addr[26531]= 1234876957;
assign addr[26532]= 1171527280;
assign addr[26533]= 1106691431;
assign addr[26534]= 1040451659;
assign addr[26535]= 972891995;
assign addr[26536]= 904098143;
assign addr[26537]= 834157373;
assign addr[26538]= 763158411;
assign addr[26539]= 691191324;
assign addr[26540]= 618347408;
assign addr[26541]= 544719071;
assign addr[26542]= 470399716;
assign addr[26543]= 395483624;
assign addr[26544]= 320065829;
assign addr[26545]= 244242007;
assign addr[26546]= 168108346;
assign addr[26547]= 91761426;
assign addr[26548]= 15298099;
assign addr[26549]= -61184634;
assign addr[26550]= -137589750;
assign addr[26551]= -213820322;
assign addr[26552]= -289779648;
assign addr[26553]= -365371365;
assign addr[26554]= -440499581;
assign addr[26555]= -515068990;
assign addr[26556]= -588984994;
assign addr[26557]= -662153826;
assign addr[26558]= -734482665;
assign addr[26559]= -805879757;
assign addr[26560]= -876254528;
assign addr[26561]= -945517704;
assign addr[26562]= -1013581418;
assign addr[26563]= -1080359326;
assign addr[26564]= -1145766716;
assign addr[26565]= -1209720613;
assign addr[26566]= -1272139887;
assign addr[26567]= -1332945355;
assign addr[26568]= -1392059879;
assign addr[26569]= -1449408469;
assign addr[26570]= -1504918373;
assign addr[26571]= -1558519173;
assign addr[26572]= -1610142873;
assign addr[26573]= -1659723983;
assign addr[26574]= -1707199606;
assign addr[26575]= -1752509516;
assign addr[26576]= -1795596234;
assign addr[26577]= -1836405100;
assign addr[26578]= -1874884346;
assign addr[26579]= -1910985158;
assign addr[26580]= -1944661739;
assign addr[26581]= -1975871368;
assign addr[26582]= -2004574453;
assign addr[26583]= -2030734582;
assign addr[26584]= -2054318569;
assign addr[26585]= -2075296495;
assign addr[26586]= -2093641749;
assign addr[26587]= -2109331059;
assign addr[26588]= -2122344521;
assign addr[26589]= -2132665626;
assign addr[26590]= -2140281282;
assign addr[26591]= -2145181827;
assign addr[26592]= -2147361045;
assign addr[26593]= -2146816171;
assign addr[26594]= -2143547897;
assign addr[26595]= -2137560369;
assign addr[26596]= -2128861181;
assign addr[26597]= -2117461370;
assign addr[26598]= -2103375398;
assign addr[26599]= -2086621133;
assign addr[26600]= -2067219829;
assign addr[26601]= -2045196100;
assign addr[26602]= -2020577882;
assign addr[26603]= -1993396407;
assign addr[26604]= -1963686155;
assign addr[26605]= -1931484818;
assign addr[26606]= -1896833245;
assign addr[26607]= -1859775393;
assign addr[26608]= -1820358275;
assign addr[26609]= -1778631892;
assign addr[26610]= -1734649179;
assign addr[26611]= -1688465931;
assign addr[26612]= -1640140734;
assign addr[26613]= -1589734894;
assign addr[26614]= -1537312353;
assign addr[26615]= -1482939614;
assign addr[26616]= -1426685652;
assign addr[26617]= -1368621831;
assign addr[26618]= -1308821808;
assign addr[26619]= -1247361445;
assign addr[26620]= -1184318708;
assign addr[26621]= -1119773573;
assign addr[26622]= -1053807919;
assign addr[26623]= -986505429;
assign addr[26624]= -917951481;
assign addr[26625]= -848233042;
assign addr[26626]= -777438554;
assign addr[26627]= -705657826;
assign addr[26628]= -632981917;
assign addr[26629]= -559503022;
assign addr[26630]= -485314355;
assign addr[26631]= -410510029;
assign addr[26632]= -335184940;
assign addr[26633]= -259434643;
assign addr[26634]= -183355234;
assign addr[26635]= -107043224;
assign addr[26636]= -30595422;
assign addr[26637]= 45891193;
assign addr[26638]= 122319591;
assign addr[26639]= 198592817;
assign addr[26640]= 274614114;
assign addr[26641]= 350287041;
assign addr[26642]= 425515602;
assign addr[26643]= 500204365;
assign addr[26644]= 574258580;
assign addr[26645]= 647584304;
assign addr[26646]= 720088517;
assign addr[26647]= 791679244;
assign addr[26648]= 862265664;
assign addr[26649]= 931758235;
assign addr[26650]= 1000068799;
assign addr[26651]= 1067110699;
assign addr[26652]= 1132798888;
assign addr[26653]= 1197050035;
assign addr[26654]= 1259782632;
assign addr[26655]= 1320917099;
assign addr[26656]= 1380375881;
assign addr[26657]= 1438083551;
assign addr[26658]= 1493966902;
assign addr[26659]= 1547955041;
assign addr[26660]= 1599979481;
assign addr[26661]= 1649974225;
assign addr[26662]= 1697875851;
assign addr[26663]= 1743623590;
assign addr[26664]= 1787159411;
assign addr[26665]= 1828428082;
assign addr[26666]= 1867377253;
assign addr[26667]= 1903957513;
assign addr[26668]= 1938122457;
assign addr[26669]= 1969828744;
assign addr[26670]= 1999036154;
assign addr[26671]= 2025707632;
assign addr[26672]= 2049809346;
assign addr[26673]= 2071310720;
assign addr[26674]= 2090184478;
assign addr[26675]= 2106406677;
assign addr[26676]= 2119956737;
assign addr[26677]= 2130817471;
assign addr[26678]= 2138975100;
assign addr[26679]= 2144419275;
assign addr[26680]= 2147143090;
assign addr[26681]= 2147143090;
assign addr[26682]= 2144419275;
assign addr[26683]= 2138975100;
assign addr[26684]= 2130817471;
assign addr[26685]= 2119956737;
assign addr[26686]= 2106406677;
assign addr[26687]= 2090184478;
assign addr[26688]= 2071310720;
assign addr[26689]= 2049809346;
assign addr[26690]= 2025707632;
assign addr[26691]= 1999036154;
assign addr[26692]= 1969828744;
assign addr[26693]= 1938122457;
assign addr[26694]= 1903957513;
assign addr[26695]= 1867377253;
assign addr[26696]= 1828428082;
assign addr[26697]= 1787159411;
assign addr[26698]= 1743623590;
assign addr[26699]= 1697875851;
assign addr[26700]= 1649974225;
assign addr[26701]= 1599979481;
assign addr[26702]= 1547955041;
assign addr[26703]= 1493966902;
assign addr[26704]= 1438083551;
assign addr[26705]= 1380375881;
assign addr[26706]= 1320917099;
assign addr[26707]= 1259782632;
assign addr[26708]= 1197050035;
assign addr[26709]= 1132798888;
assign addr[26710]= 1067110699;
assign addr[26711]= 1000068799;
assign addr[26712]= 931758235;
assign addr[26713]= 862265664;
assign addr[26714]= 791679244;
assign addr[26715]= 720088517;
assign addr[26716]= 647584304;
assign addr[26717]= 574258580;
assign addr[26718]= 500204365;
assign addr[26719]= 425515602;
assign addr[26720]= 350287041;
assign addr[26721]= 274614114;
assign addr[26722]= 198592817;
assign addr[26723]= 122319591;
assign addr[26724]= 45891193;
assign addr[26725]= -30595422;
assign addr[26726]= -107043224;
assign addr[26727]= -183355234;
assign addr[26728]= -259434643;
assign addr[26729]= -335184940;
assign addr[26730]= -410510029;
assign addr[26731]= -485314355;
assign addr[26732]= -559503022;
assign addr[26733]= -632981917;
assign addr[26734]= -705657826;
assign addr[26735]= -777438554;
assign addr[26736]= -848233042;
assign addr[26737]= -917951481;
assign addr[26738]= -986505429;
assign addr[26739]= -1053807919;
assign addr[26740]= -1119773573;
assign addr[26741]= -1184318708;
assign addr[26742]= -1247361445;
assign addr[26743]= -1308821808;
assign addr[26744]= -1368621831;
assign addr[26745]= -1426685652;
assign addr[26746]= -1482939614;
assign addr[26747]= -1537312353;
assign addr[26748]= -1589734894;
assign addr[26749]= -1640140734;
assign addr[26750]= -1688465931;
assign addr[26751]= -1734649179;
assign addr[26752]= -1778631892;
assign addr[26753]= -1820358275;
assign addr[26754]= -1859775393;
assign addr[26755]= -1896833245;
assign addr[26756]= -1931484818;
assign addr[26757]= -1963686155;
assign addr[26758]= -1993396407;
assign addr[26759]= -2020577882;
assign addr[26760]= -2045196100;
assign addr[26761]= -2067219829;
assign addr[26762]= -2086621133;
assign addr[26763]= -2103375398;
assign addr[26764]= -2117461370;
assign addr[26765]= -2128861181;
assign addr[26766]= -2137560369;
assign addr[26767]= -2143547897;
assign addr[26768]= -2146816171;
assign addr[26769]= -2147361045;
assign addr[26770]= -2145181827;
assign addr[26771]= -2140281282;
assign addr[26772]= -2132665626;
assign addr[26773]= -2122344521;
assign addr[26774]= -2109331059;
assign addr[26775]= -2093641749;
assign addr[26776]= -2075296495;
assign addr[26777]= -2054318569;
assign addr[26778]= -2030734582;
assign addr[26779]= -2004574453;
assign addr[26780]= -1975871368;
assign addr[26781]= -1944661739;
assign addr[26782]= -1910985158;
assign addr[26783]= -1874884346;
assign addr[26784]= -1836405100;
assign addr[26785]= -1795596234;
assign addr[26786]= -1752509516;
assign addr[26787]= -1707199606;
assign addr[26788]= -1659723983;
assign addr[26789]= -1610142873;
assign addr[26790]= -1558519173;
assign addr[26791]= -1504918373;
assign addr[26792]= -1449408469;
assign addr[26793]= -1392059879;
assign addr[26794]= -1332945355;
assign addr[26795]= -1272139887;
assign addr[26796]= -1209720613;
assign addr[26797]= -1145766716;
assign addr[26798]= -1080359326;
assign addr[26799]= -1013581418;
assign addr[26800]= -945517704;
assign addr[26801]= -876254528;
assign addr[26802]= -805879757;
assign addr[26803]= -734482665;
assign addr[26804]= -662153826;
assign addr[26805]= -588984994;
assign addr[26806]= -515068990;
assign addr[26807]= -440499581;
assign addr[26808]= -365371365;
assign addr[26809]= -289779648;
assign addr[26810]= -213820322;
assign addr[26811]= -137589750;
assign addr[26812]= -61184634;
assign addr[26813]= 15298099;
assign addr[26814]= 91761426;
assign addr[26815]= 168108346;
assign addr[26816]= 244242007;
assign addr[26817]= 320065829;
assign addr[26818]= 395483624;
assign addr[26819]= 470399716;
assign addr[26820]= 544719071;
assign addr[26821]= 618347408;
assign addr[26822]= 691191324;
assign addr[26823]= 763158411;
assign addr[26824]= 834157373;
assign addr[26825]= 904098143;
assign addr[26826]= 972891995;
assign addr[26827]= 1040451659;
assign addr[26828]= 1106691431;
assign addr[26829]= 1171527280;
assign addr[26830]= 1234876957;
assign addr[26831]= 1296660098;
assign addr[26832]= 1356798326;
assign addr[26833]= 1415215352;
assign addr[26834]= 1471837070;
assign addr[26835]= 1526591649;
assign addr[26836]= 1579409630;
assign addr[26837]= 1630224009;
assign addr[26838]= 1678970324;
assign addr[26839]= 1725586737;
assign addr[26840]= 1770014111;
assign addr[26841]= 1812196087;
assign addr[26842]= 1852079154;
assign addr[26843]= 1889612716;
assign addr[26844]= 1924749160;
assign addr[26845]= 1957443913;
assign addr[26846]= 1987655498;
assign addr[26847]= 2015345591;
assign addr[26848]= 2040479063;
assign addr[26849]= 2063024031;
assign addr[26850]= 2082951896;
assign addr[26851]= 2100237377;
assign addr[26852]= 2114858546;
assign addr[26853]= 2126796855;
assign addr[26854]= 2136037160;
assign addr[26855]= 2142567738;
assign addr[26856]= 2146380306;
assign addr[26857]= 2147470025;
assign addr[26858]= 2145835515;
assign addr[26859]= 2141478848;
assign addr[26860]= 2134405552;
assign addr[26861]= 2124624598;
assign addr[26862]= 2112148396;
assign addr[26863]= 2096992772;
assign addr[26864]= 2079176953;
assign addr[26865]= 2058723538;
assign addr[26866]= 2035658475;
assign addr[26867]= 2010011024;
assign addr[26868]= 1981813720;
assign addr[26869]= 1951102334;
assign addr[26870]= 1917915825;
assign addr[26871]= 1882296293;
assign addr[26872]= 1844288924;
assign addr[26873]= 1803941934;
assign addr[26874]= 1761306505;
assign addr[26875]= 1716436725;
assign addr[26876]= 1669389513;
assign addr[26877]= 1620224553;
assign addr[26878]= 1569004214;
assign addr[26879]= 1515793473;
assign addr[26880]= 1460659832;
assign addr[26881]= 1403673233;
assign addr[26882]= 1344905966;
assign addr[26883]= 1284432584;
assign addr[26884]= 1222329801;
assign addr[26885]= 1158676398;
assign addr[26886]= 1093553126;
assign addr[26887]= 1027042599;
assign addr[26888]= 959229189;
assign addr[26889]= 890198924;
assign addr[26890]= 820039373;
assign addr[26891]= 748839539;
assign addr[26892]= 676689746;
assign addr[26893]= 603681519;
assign addr[26894]= 529907477;
assign addr[26895]= 455461206;
assign addr[26896]= 380437148;
assign addr[26897]= 304930476;
assign addr[26898]= 229036977;
assign addr[26899]= 152852926;
assign addr[26900]= 76474970;
assign addr[26901]= 0;
assign addr[26902]= -76474970;
assign addr[26903]= -152852926;
assign addr[26904]= -229036977;
assign addr[26905]= -304930476;
assign addr[26906]= -380437148;
assign addr[26907]= -455461206;
assign addr[26908]= -529907477;
assign addr[26909]= -603681519;
assign addr[26910]= -676689746;
assign addr[26911]= -748839539;
assign addr[26912]= -820039373;
assign addr[26913]= -890198924;
assign addr[26914]= -959229189;
assign addr[26915]= -1027042599;
assign addr[26916]= -1093553126;
assign addr[26917]= -1158676398;
assign addr[26918]= -1222329801;
assign addr[26919]= -1284432584;
assign addr[26920]= -1344905966;
assign addr[26921]= -1403673233;
assign addr[26922]= -1460659832;
assign addr[26923]= -1515793473;
assign addr[26924]= -1569004214;
assign addr[26925]= -1620224553;
assign addr[26926]= -1669389513;
assign addr[26927]= -1716436725;
assign addr[26928]= -1761306505;
assign addr[26929]= -1803941934;
assign addr[26930]= -1844288924;
assign addr[26931]= -1882296293;
assign addr[26932]= -1917915825;
assign addr[26933]= -1951102334;
assign addr[26934]= -1981813720;
assign addr[26935]= -2010011024;
assign addr[26936]= -2035658475;
assign addr[26937]= -2058723538;
assign addr[26938]= -2079176953;
assign addr[26939]= -2096992772;
assign addr[26940]= -2112148396;
assign addr[26941]= -2124624598;
assign addr[26942]= -2134405552;
assign addr[26943]= -2141478848;
assign addr[26944]= -2145835515;
assign addr[26945]= -2147470025;
assign addr[26946]= -2146380306;
assign addr[26947]= -2142567738;
assign addr[26948]= -2136037160;
assign addr[26949]= -2126796855;
assign addr[26950]= -2114858546;
assign addr[26951]= -2100237377;
assign addr[26952]= -2082951896;
assign addr[26953]= -2063024031;
assign addr[26954]= -2040479063;
assign addr[26955]= -2015345591;
assign addr[26956]= -1987655498;
assign addr[26957]= -1957443913;
assign addr[26958]= -1924749160;
assign addr[26959]= -1889612716;
assign addr[26960]= -1852079154;
assign addr[26961]= -1812196087;
assign addr[26962]= -1770014111;
assign addr[26963]= -1725586737;
assign addr[26964]= -1678970324;
assign addr[26965]= -1630224009;
assign addr[26966]= -1579409630;
assign addr[26967]= -1526591649;
assign addr[26968]= -1471837070;
assign addr[26969]= -1415215352;
assign addr[26970]= -1356798326;
assign addr[26971]= -1296660098;
assign addr[26972]= -1234876957;
assign addr[26973]= -1171527280;
assign addr[26974]= -1106691431;
assign addr[26975]= -1040451659;
assign addr[26976]= -972891995;
assign addr[26977]= -904098143;
assign addr[26978]= -834157373;
assign addr[26979]= -763158411;
assign addr[26980]= -691191324;
assign addr[26981]= -618347408;
assign addr[26982]= -544719071;
assign addr[26983]= -470399716;
assign addr[26984]= -395483624;
assign addr[26985]= -320065829;
assign addr[26986]= -244242007;
assign addr[26987]= -168108346;
assign addr[26988]= -91761426;
assign addr[26989]= -15298099;
assign addr[26990]= 61184634;
assign addr[26991]= 137589750;
assign addr[26992]= 213820322;
assign addr[26993]= 289779648;
assign addr[26994]= 365371365;
assign addr[26995]= 440499581;
assign addr[26996]= 515068990;
assign addr[26997]= 588984994;
assign addr[26998]= 662153826;
assign addr[26999]= 734482665;
assign addr[27000]= 805879757;
assign addr[27001]= 876254528;
assign addr[27002]= 945517704;
assign addr[27003]= 1013581418;
assign addr[27004]= 1080359326;
assign addr[27005]= 1145766716;
assign addr[27006]= 1209720613;
assign addr[27007]= 1272139887;
assign addr[27008]= 1332945355;
assign addr[27009]= 1392059879;
assign addr[27010]= 1449408469;
assign addr[27011]= 1504918373;
assign addr[27012]= 1558519173;
assign addr[27013]= 1610142873;
assign addr[27014]= 1659723983;
assign addr[27015]= 1707199606;
assign addr[27016]= 1752509516;
assign addr[27017]= 1795596234;
assign addr[27018]= 1836405100;
assign addr[27019]= 1874884346;
assign addr[27020]= 1910985158;
assign addr[27021]= 1944661739;
assign addr[27022]= 1975871368;
assign addr[27023]= 2004574453;
assign addr[27024]= 2030734582;
assign addr[27025]= 2054318569;
assign addr[27026]= 2075296495;
assign addr[27027]= 2093641749;
assign addr[27028]= 2109331059;
assign addr[27029]= 2122344521;
assign addr[27030]= 2132665626;
assign addr[27031]= 2140281282;
assign addr[27032]= 2145181827;
assign addr[27033]= 2147361045;
assign addr[27034]= 2146816171;
assign addr[27035]= 2143547897;
assign addr[27036]= 2137560369;
assign addr[27037]= 2128861181;
assign addr[27038]= 2117461370;
assign addr[27039]= 2103375398;
assign addr[27040]= 2086621133;
assign addr[27041]= 2067219829;
assign addr[27042]= 2045196100;
assign addr[27043]= 2020577882;
assign addr[27044]= 1993396407;
assign addr[27045]= 1963686155;
assign addr[27046]= 1931484818;
assign addr[27047]= 1896833245;
assign addr[27048]= 1859775393;
assign addr[27049]= 1820358275;
assign addr[27050]= 1778631892;
assign addr[27051]= 1734649179;
assign addr[27052]= 1688465931;
assign addr[27053]= 1640140734;
assign addr[27054]= 1589734894;
assign addr[27055]= 1537312353;
assign addr[27056]= 1482939614;
assign addr[27057]= 1426685652;
assign addr[27058]= 1368621831;
assign addr[27059]= 1308821808;
assign addr[27060]= 1247361445;
assign addr[27061]= 1184318708;
assign addr[27062]= 1119773573;
assign addr[27063]= 1053807919;
assign addr[27064]= 986505429;
assign addr[27065]= 917951481;
assign addr[27066]= 848233042;
assign addr[27067]= 777438554;
assign addr[27068]= 705657826;
assign addr[27069]= 632981917;
assign addr[27070]= 559503022;
assign addr[27071]= 485314355;
assign addr[27072]= 410510029;
assign addr[27073]= 335184940;
assign addr[27074]= 259434643;
assign addr[27075]= 183355234;
assign addr[27076]= 107043224;
assign addr[27077]= 30595422;
assign addr[27078]= -45891193;
assign addr[27079]= -122319591;
assign addr[27080]= -198592817;
assign addr[27081]= -274614114;
assign addr[27082]= -350287041;
assign addr[27083]= -425515602;
assign addr[27084]= -500204365;
assign addr[27085]= -574258580;
assign addr[27086]= -647584304;
assign addr[27087]= -720088517;
assign addr[27088]= -791679244;
assign addr[27089]= -862265664;
assign addr[27090]= -931758235;
assign addr[27091]= -1000068799;
assign addr[27092]= -1067110699;
assign addr[27093]= -1132798888;
assign addr[27094]= -1197050035;
assign addr[27095]= -1259782632;
assign addr[27096]= -1320917099;
assign addr[27097]= -1380375881;
assign addr[27098]= -1438083551;
assign addr[27099]= -1493966902;
assign addr[27100]= -1547955041;
assign addr[27101]= -1599979481;
assign addr[27102]= -1649974225;
assign addr[27103]= -1697875851;
assign addr[27104]= -1743623590;
assign addr[27105]= -1787159411;
assign addr[27106]= -1828428082;
assign addr[27107]= -1867377253;
assign addr[27108]= -1903957513;
assign addr[27109]= -1938122457;
assign addr[27110]= -1969828744;
assign addr[27111]= -1999036154;
assign addr[27112]= -2025707632;
assign addr[27113]= -2049809346;
assign addr[27114]= -2071310720;
assign addr[27115]= -2090184478;
assign addr[27116]= -2106406677;
assign addr[27117]= -2119956737;
assign addr[27118]= -2130817471;
assign addr[27119]= -2138975100;
assign addr[27120]= -2144419275;
assign addr[27121]= -2147143090;
assign addr[27122]= -2147143090;
assign addr[27123]= -2144419275;
assign addr[27124]= -2138975100;
assign addr[27125]= -2130817471;
assign addr[27126]= -2119956737;
assign addr[27127]= -2106406677;
assign addr[27128]= -2090184478;
assign addr[27129]= -2071310720;
assign addr[27130]= -2049809346;
assign addr[27131]= -2025707632;
assign addr[27132]= -1999036154;
assign addr[27133]= -1969828744;
assign addr[27134]= -1938122457;
assign addr[27135]= -1903957513;
assign addr[27136]= -1867377253;
assign addr[27137]= -1828428082;
assign addr[27138]= -1787159411;
assign addr[27139]= -1743623590;
assign addr[27140]= -1697875851;
assign addr[27141]= -1649974225;
assign addr[27142]= -1599979481;
assign addr[27143]= -1547955041;
assign addr[27144]= -1493966902;
assign addr[27145]= -1438083551;
assign addr[27146]= -1380375881;
assign addr[27147]= -1320917099;
assign addr[27148]= -1259782632;
assign addr[27149]= -1197050035;
assign addr[27150]= -1132798888;
assign addr[27151]= -1067110699;
assign addr[27152]= -1000068799;
assign addr[27153]= -931758235;
assign addr[27154]= -862265664;
assign addr[27155]= -791679244;
assign addr[27156]= -720088517;
assign addr[27157]= -647584304;
assign addr[27158]= -574258580;
assign addr[27159]= -500204365;
assign addr[27160]= -425515602;
assign addr[27161]= -350287041;
assign addr[27162]= -274614114;
assign addr[27163]= -198592817;
assign addr[27164]= -122319591;
assign addr[27165]= -45891193;
assign addr[27166]= 30595422;
assign addr[27167]= 107043224;
assign addr[27168]= 183355234;
assign addr[27169]= 259434643;
assign addr[27170]= 335184940;
assign addr[27171]= 410510029;
assign addr[27172]= 485314355;
assign addr[27173]= 559503022;
assign addr[27174]= 632981917;
assign addr[27175]= 705657826;
assign addr[27176]= 777438554;
assign addr[27177]= 848233042;
assign addr[27178]= 917951481;
assign addr[27179]= 986505429;
assign addr[27180]= 1053807919;
assign addr[27181]= 1119773573;
assign addr[27182]= 1184318708;
assign addr[27183]= 1247361445;
assign addr[27184]= 1308821808;
assign addr[27185]= 1368621831;
assign addr[27186]= 1426685652;
assign addr[27187]= 1482939614;
assign addr[27188]= 1537312353;
assign addr[27189]= 1589734894;
assign addr[27190]= 1640140734;
assign addr[27191]= 1688465931;
assign addr[27192]= 1734649179;
assign addr[27193]= 1778631892;
assign addr[27194]= 1820358275;
assign addr[27195]= 1859775393;
assign addr[27196]= 1896833245;
assign addr[27197]= 1931484818;
assign addr[27198]= 1963686155;
assign addr[27199]= 1993396407;
assign addr[27200]= 2020577882;
assign addr[27201]= 2045196100;
assign addr[27202]= 2067219829;
assign addr[27203]= 2086621133;
assign addr[27204]= 2103375398;
assign addr[27205]= 2117461370;
assign addr[27206]= 2128861181;
assign addr[27207]= 2137560369;
assign addr[27208]= 2143547897;
assign addr[27209]= 2146816171;
assign addr[27210]= 2147361045;
assign addr[27211]= 2145181827;
assign addr[27212]= 2140281282;
assign addr[27213]= 2132665626;
assign addr[27214]= 2122344521;
assign addr[27215]= 2109331059;
assign addr[27216]= 2093641749;
assign addr[27217]= 2075296495;
assign addr[27218]= 2054318569;
assign addr[27219]= 2030734582;
assign addr[27220]= 2004574453;
assign addr[27221]= 1975871368;
assign addr[27222]= 1944661739;
assign addr[27223]= 1910985158;
assign addr[27224]= 1874884346;
assign addr[27225]= 1836405100;
assign addr[27226]= 1795596234;
assign addr[27227]= 1752509516;
assign addr[27228]= 1707199606;
assign addr[27229]= 1659723983;
assign addr[27230]= 1610142873;
assign addr[27231]= 1558519173;
assign addr[27232]= 1504918373;
assign addr[27233]= 1449408469;
assign addr[27234]= 1392059879;
assign addr[27235]= 1332945355;
assign addr[27236]= 1272139887;
assign addr[27237]= 1209720613;
assign addr[27238]= 1145766716;
assign addr[27239]= 1080359326;
assign addr[27240]= 1013581418;
assign addr[27241]= 945517704;
assign addr[27242]= 876254528;
assign addr[27243]= 805879757;
assign addr[27244]= 734482665;
assign addr[27245]= 662153826;
assign addr[27246]= 588984994;
assign addr[27247]= 515068990;
assign addr[27248]= 440499581;
assign addr[27249]= 365371365;
assign addr[27250]= 289779648;
assign addr[27251]= 213820322;
assign addr[27252]= 137589750;
assign addr[27253]= 61184634;
assign addr[27254]= -15298099;
assign addr[27255]= -91761426;
assign addr[27256]= -168108346;
assign addr[27257]= -244242007;
assign addr[27258]= -320065829;
assign addr[27259]= -395483624;
assign addr[27260]= -470399716;
assign addr[27261]= -544719071;
assign addr[27262]= -618347408;
assign addr[27263]= -691191324;
assign addr[27264]= -763158411;
assign addr[27265]= -834157373;
assign addr[27266]= -904098143;
assign addr[27267]= -972891995;
assign addr[27268]= -1040451659;
assign addr[27269]= -1106691431;
assign addr[27270]= -1171527280;
assign addr[27271]= -1234876957;
assign addr[27272]= -1296660098;
assign addr[27273]= -1356798326;
assign addr[27274]= -1415215352;
assign addr[27275]= -1471837070;
assign addr[27276]= -1526591649;
assign addr[27277]= -1579409630;
assign addr[27278]= -1630224009;
assign addr[27279]= -1678970324;
assign addr[27280]= -1725586737;
assign addr[27281]= -1770014111;
assign addr[27282]= -1812196087;
assign addr[27283]= -1852079154;
assign addr[27284]= -1889612716;
assign addr[27285]= -1924749160;
assign addr[27286]= -1957443913;
assign addr[27287]= -1987655498;
assign addr[27288]= -2015345591;
assign addr[27289]= -2040479063;
assign addr[27290]= -2063024031;
assign addr[27291]= -2082951896;
assign addr[27292]= -2100237377;
assign addr[27293]= -2114858546;
assign addr[27294]= -2126796855;
assign addr[27295]= -2136037160;
assign addr[27296]= -2142567738;
assign addr[27297]= -2146380306;
assign addr[27298]= -2147470025;
assign addr[27299]= -2145835515;
assign addr[27300]= -2141478848;
assign addr[27301]= -2134405552;
assign addr[27302]= -2124624598;
assign addr[27303]= -2112148396;
assign addr[27304]= -2096992772;
assign addr[27305]= -2079176953;
assign addr[27306]= -2058723538;
assign addr[27307]= -2035658475;
assign addr[27308]= -2010011024;
assign addr[27309]= -1981813720;
assign addr[27310]= -1951102334;
assign addr[27311]= -1917915825;
assign addr[27312]= -1882296293;
assign addr[27313]= -1844288924;
assign addr[27314]= -1803941934;
assign addr[27315]= -1761306505;
assign addr[27316]= -1716436725;
assign addr[27317]= -1669389513;
assign addr[27318]= -1620224553;
assign addr[27319]= -1569004214;
assign addr[27320]= -1515793473;
assign addr[27321]= -1460659832;
assign addr[27322]= -1403673233;
assign addr[27323]= -1344905966;
assign addr[27324]= -1284432584;
assign addr[27325]= -1222329801;
assign addr[27326]= -1158676398;
assign addr[27327]= -1093553126;
assign addr[27328]= -1027042599;
assign addr[27329]= -959229189;
assign addr[27330]= -890198924;
assign addr[27331]= -820039373;
assign addr[27332]= -748839539;
assign addr[27333]= -676689746;
assign addr[27334]= -603681519;
assign addr[27335]= -529907477;
assign addr[27336]= -455461206;
assign addr[27337]= -380437148;
assign addr[27338]= -304930476;
assign addr[27339]= -229036977;
assign addr[27340]= -152852926;
assign addr[27341]= -76474970;
assign addr[27342]= 0;
assign addr[27343]= 76474970;
assign addr[27344]= 152852926;
assign addr[27345]= 229036977;
assign addr[27346]= 304930476;
assign addr[27347]= 380437148;
assign addr[27348]= 455461206;
assign addr[27349]= 529907477;
assign addr[27350]= 603681519;
assign addr[27351]= 676689746;
assign addr[27352]= 748839539;
assign addr[27353]= 820039373;
assign addr[27354]= 890198924;
assign addr[27355]= 959229189;
assign addr[27356]= 1027042599;
assign addr[27357]= 1093553126;
assign addr[27358]= 1158676398;
assign addr[27359]= 1222329801;
assign addr[27360]= 1284432584;
assign addr[27361]= 1344905966;
assign addr[27362]= 1403673233;
assign addr[27363]= 1460659832;
assign addr[27364]= 1515793473;
assign addr[27365]= 1569004214;
assign addr[27366]= 1620224553;
assign addr[27367]= 1669389513;
assign addr[27368]= 1716436725;
assign addr[27369]= 1761306505;
assign addr[27370]= 1803941934;
assign addr[27371]= 1844288924;
assign addr[27372]= 1882296293;
assign addr[27373]= 1917915825;
assign addr[27374]= 1951102334;
assign addr[27375]= 1981813720;
assign addr[27376]= 2010011024;
assign addr[27377]= 2035658475;
assign addr[27378]= 2058723538;
assign addr[27379]= 2079176953;
assign addr[27380]= 2096992772;
assign addr[27381]= 2112148396;
assign addr[27382]= 2124624598;
assign addr[27383]= 2134405552;
assign addr[27384]= 2141478848;
assign addr[27385]= 2145835515;
assign addr[27386]= 2147470025;
assign addr[27387]= 2146380306;
assign addr[27388]= 2142567738;
assign addr[27389]= 2136037160;
assign addr[27390]= 2126796855;
assign addr[27391]= 2114858546;
assign addr[27392]= 2100237377;
assign addr[27393]= 2082951896;
assign addr[27394]= 2063024031;
assign addr[27395]= 2040479063;
assign addr[27396]= 2015345591;
assign addr[27397]= 1987655498;
assign addr[27398]= 1957443913;
assign addr[27399]= 1924749160;
assign addr[27400]= 1889612716;
assign addr[27401]= 1852079154;
assign addr[27402]= 1812196087;
assign addr[27403]= 1770014111;
assign addr[27404]= 1725586737;
assign addr[27405]= 1678970324;
assign addr[27406]= 1630224009;
assign addr[27407]= 1579409630;
assign addr[27408]= 1526591649;
assign addr[27409]= 1471837070;
assign addr[27410]= 1415215352;
assign addr[27411]= 1356798326;
assign addr[27412]= 1296660098;
assign addr[27413]= 1234876957;
assign addr[27414]= 1171527280;
assign addr[27415]= 1106691431;
assign addr[27416]= 1040451659;
assign addr[27417]= 972891995;
assign addr[27418]= 904098143;
assign addr[27419]= 834157373;
assign addr[27420]= 763158411;
assign addr[27421]= 691191324;
assign addr[27422]= 618347408;
assign addr[27423]= 544719071;
assign addr[27424]= 470399716;
assign addr[27425]= 395483624;
assign addr[27426]= 320065829;
assign addr[27427]= 244242007;
assign addr[27428]= 168108346;
assign addr[27429]= 91761426;
assign addr[27430]= 15298099;
assign addr[27431]= -61184634;
assign addr[27432]= -137589750;
assign addr[27433]= -213820322;
assign addr[27434]= -289779648;
assign addr[27435]= -365371365;
assign addr[27436]= -440499581;
assign addr[27437]= -515068990;
assign addr[27438]= -588984994;
assign addr[27439]= -662153826;
assign addr[27440]= -734482665;
assign addr[27441]= -805879757;
assign addr[27442]= -876254528;
assign addr[27443]= -945517704;
assign addr[27444]= -1013581418;
assign addr[27445]= -1080359326;
assign addr[27446]= -1145766716;
assign addr[27447]= -1209720613;
assign addr[27448]= -1272139887;
assign addr[27449]= -1332945355;
assign addr[27450]= -1392059879;
assign addr[27451]= -1449408469;
assign addr[27452]= -1504918373;
assign addr[27453]= -1558519173;
assign addr[27454]= -1610142873;
assign addr[27455]= -1659723983;
assign addr[27456]= -1707199606;
assign addr[27457]= -1752509516;
assign addr[27458]= -1795596234;
assign addr[27459]= -1836405100;
assign addr[27460]= -1874884346;
assign addr[27461]= -1910985158;
assign addr[27462]= -1944661739;
assign addr[27463]= -1975871368;
assign addr[27464]= -2004574453;
assign addr[27465]= -2030734582;
assign addr[27466]= -2054318569;
assign addr[27467]= -2075296495;
assign addr[27468]= -2093641749;
assign addr[27469]= -2109331059;
assign addr[27470]= -2122344521;
assign addr[27471]= -2132665626;
assign addr[27472]= -2140281282;
assign addr[27473]= -2145181827;
assign addr[27474]= -2147361045;
assign addr[27475]= -2146816171;
assign addr[27476]= -2143547897;
assign addr[27477]= -2137560369;
assign addr[27478]= -2128861181;
assign addr[27479]= -2117461370;
assign addr[27480]= -2103375398;
assign addr[27481]= -2086621133;
assign addr[27482]= -2067219829;
assign addr[27483]= -2045196100;
assign addr[27484]= -2020577882;
assign addr[27485]= -1993396407;
assign addr[27486]= -1963686155;
assign addr[27487]= -1931484818;
assign addr[27488]= -1896833245;
assign addr[27489]= -1859775393;
assign addr[27490]= -1820358275;
assign addr[27491]= -1778631892;
assign addr[27492]= -1734649179;
assign addr[27493]= -1688465931;
assign addr[27494]= -1640140734;
assign addr[27495]= -1589734894;
assign addr[27496]= -1537312353;
assign addr[27497]= -1482939614;
assign addr[27498]= -1426685652;
assign addr[27499]= -1368621831;
assign addr[27500]= -1308821808;
assign addr[27501]= -1247361445;
assign addr[27502]= -1184318708;
assign addr[27503]= -1119773573;
assign addr[27504]= -1053807919;
assign addr[27505]= -986505429;
assign addr[27506]= -917951481;
assign addr[27507]= -848233042;
assign addr[27508]= -777438554;
assign addr[27509]= -705657826;
assign addr[27510]= -632981917;
assign addr[27511]= -559503022;
assign addr[27512]= -485314355;
assign addr[27513]= -410510029;
assign addr[27514]= -335184940;
assign addr[27515]= -259434643;
assign addr[27516]= -183355234;
assign addr[27517]= -107043224;
assign addr[27518]= -30595422;
assign addr[27519]= 45891193;
assign addr[27520]= 122319591;
assign addr[27521]= 198592817;
assign addr[27522]= 274614114;
assign addr[27523]= 350287041;
assign addr[27524]= 425515602;
assign addr[27525]= 500204365;
assign addr[27526]= 574258580;
assign addr[27527]= 647584304;
assign addr[27528]= 720088517;
assign addr[27529]= 791679244;
assign addr[27530]= 862265664;
assign addr[27531]= 931758235;
assign addr[27532]= 1000068799;
assign addr[27533]= 1067110699;
assign addr[27534]= 1132798888;
assign addr[27535]= 1197050035;
assign addr[27536]= 1259782632;
assign addr[27537]= 1320917099;
assign addr[27538]= 1380375881;
assign addr[27539]= 1438083551;
assign addr[27540]= 1493966902;
assign addr[27541]= 1547955041;
assign addr[27542]= 1599979481;
assign addr[27543]= 1649974225;
assign addr[27544]= 1697875851;
assign addr[27545]= 1743623590;
assign addr[27546]= 1787159411;
assign addr[27547]= 1828428082;
assign addr[27548]= 1867377253;
assign addr[27549]= 1903957513;
assign addr[27550]= 1938122457;
assign addr[27551]= 1969828744;
assign addr[27552]= 1999036154;
assign addr[27553]= 2025707632;
assign addr[27554]= 2049809346;
assign addr[27555]= 2071310720;
assign addr[27556]= 2090184478;
assign addr[27557]= 2106406677;
assign addr[27558]= 2119956737;
assign addr[27559]= 2130817471;
assign addr[27560]= 2138975100;
assign addr[27561]= 2144419275;
assign addr[27562]= 2147143090;
assign addr[27563]= 2147143090;
assign addr[27564]= 2144419275;
assign addr[27565]= 2138975100;
assign addr[27566]= 2130817471;
assign addr[27567]= 2119956737;
assign addr[27568]= 2106406677;
assign addr[27569]= 2090184478;
assign addr[27570]= 2071310720;
assign addr[27571]= 2049809346;
assign addr[27572]= 2025707632;
assign addr[27573]= 1999036154;
assign addr[27574]= 1969828744;
assign addr[27575]= 1938122457;
assign addr[27576]= 1903957513;
assign addr[27577]= 1867377253;
assign addr[27578]= 1828428082;
assign addr[27579]= 1787159411;
assign addr[27580]= 1743623590;
assign addr[27581]= 1697875851;
assign addr[27582]= 1649974225;
assign addr[27583]= 1599979481;
assign addr[27584]= 1547955041;
assign addr[27585]= 1493966902;
assign addr[27586]= 1438083551;
assign addr[27587]= 1380375881;
assign addr[27588]= 1320917099;
assign addr[27589]= 1259782632;
assign addr[27590]= 1197050035;
assign addr[27591]= 1132798888;
assign addr[27592]= 1067110699;
assign addr[27593]= 1000068799;
assign addr[27594]= 931758235;
assign addr[27595]= 862265664;
assign addr[27596]= 791679244;
assign addr[27597]= 720088517;
assign addr[27598]= 647584304;
assign addr[27599]= 574258580;
assign addr[27600]= 500204365;
assign addr[27601]= 425515602;
assign addr[27602]= 350287041;
assign addr[27603]= 274614114;
assign addr[27604]= 198592817;
assign addr[27605]= 122319591;
assign addr[27606]= 45891193;
assign addr[27607]= -30595422;
assign addr[27608]= -107043224;
assign addr[27609]= -183355234;
assign addr[27610]= -259434643;
assign addr[27611]= -335184940;
assign addr[27612]= -410510029;
assign addr[27613]= -485314355;
assign addr[27614]= -559503022;
assign addr[27615]= -632981917;
assign addr[27616]= -705657826;
assign addr[27617]= -777438554;
assign addr[27618]= -848233042;
assign addr[27619]= -917951481;
assign addr[27620]= -986505429;
assign addr[27621]= -1053807919;
assign addr[27622]= -1119773573;
assign addr[27623]= -1184318708;
assign addr[27624]= -1247361445;
assign addr[27625]= -1308821808;
assign addr[27626]= -1368621831;
assign addr[27627]= -1426685652;
assign addr[27628]= -1482939614;
assign addr[27629]= -1537312353;
assign addr[27630]= -1589734894;
assign addr[27631]= -1640140734;
assign addr[27632]= -1688465931;
assign addr[27633]= -1734649179;
assign addr[27634]= -1778631892;
assign addr[27635]= -1820358275;
assign addr[27636]= -1859775393;
assign addr[27637]= -1896833245;
assign addr[27638]= -1931484818;
assign addr[27639]= -1963686155;
assign addr[27640]= -1993396407;
assign addr[27641]= -2020577882;
assign addr[27642]= -2045196100;
assign addr[27643]= -2067219829;
assign addr[27644]= -2086621133;
assign addr[27645]= -2103375398;
assign addr[27646]= -2117461370;
assign addr[27647]= -2128861181;
assign addr[27648]= -2137560369;
assign addr[27649]= -2143547897;
assign addr[27650]= -2146816171;
assign addr[27651]= -2147361045;
assign addr[27652]= -2145181827;
assign addr[27653]= -2140281282;
assign addr[27654]= -2132665626;
assign addr[27655]= -2122344521;
assign addr[27656]= -2109331059;
assign addr[27657]= -2093641749;
assign addr[27658]= -2075296495;
assign addr[27659]= -2054318569;
assign addr[27660]= -2030734582;
assign addr[27661]= -2004574453;
assign addr[27662]= -1975871368;
assign addr[27663]= -1944661739;
assign addr[27664]= -1910985158;
assign addr[27665]= -1874884346;
assign addr[27666]= -1836405100;
assign addr[27667]= -1795596234;
assign addr[27668]= -1752509516;
assign addr[27669]= -1707199606;
assign addr[27670]= -1659723983;
assign addr[27671]= -1610142873;
assign addr[27672]= -1558519173;
assign addr[27673]= -1504918373;
assign addr[27674]= -1449408469;
assign addr[27675]= -1392059879;
assign addr[27676]= -1332945355;
assign addr[27677]= -1272139887;
assign addr[27678]= -1209720613;
assign addr[27679]= -1145766716;
assign addr[27680]= -1080359326;
assign addr[27681]= -1013581418;
assign addr[27682]= -945517704;
assign addr[27683]= -876254528;
assign addr[27684]= -805879757;
assign addr[27685]= -734482665;
assign addr[27686]= -662153826;
assign addr[27687]= -588984994;
assign addr[27688]= -515068990;
assign addr[27689]= -440499581;
assign addr[27690]= -365371365;
assign addr[27691]= -289779648;
assign addr[27692]= -213820322;
assign addr[27693]= -137589750;
assign addr[27694]= -61184634;
assign addr[27695]= 15298099;
assign addr[27696]= 91761426;
assign addr[27697]= 168108346;
assign addr[27698]= 244242007;
assign addr[27699]= 320065829;
assign addr[27700]= 395483624;
assign addr[27701]= 470399716;
assign addr[27702]= 544719071;
assign addr[27703]= 618347408;
assign addr[27704]= 691191324;
assign addr[27705]= 763158411;
assign addr[27706]= 834157373;
assign addr[27707]= 904098143;
assign addr[27708]= 972891995;
assign addr[27709]= 1040451659;
assign addr[27710]= 1106691431;
assign addr[27711]= 1171527280;
assign addr[27712]= 1234876957;
assign addr[27713]= 1296660098;
assign addr[27714]= 1356798326;
assign addr[27715]= 1415215352;
assign addr[27716]= 1471837070;
assign addr[27717]= 1526591649;
assign addr[27718]= 1579409630;
assign addr[27719]= 1630224009;
assign addr[27720]= 1678970324;
assign addr[27721]= 1725586737;
assign addr[27722]= 1770014111;
assign addr[27723]= 1812196087;
assign addr[27724]= 1852079154;
assign addr[27725]= 1889612716;
assign addr[27726]= 1924749160;
assign addr[27727]= 1957443913;
assign addr[27728]= 1987655498;
assign addr[27729]= 2015345591;
assign addr[27730]= 2040479063;
assign addr[27731]= 2063024031;
assign addr[27732]= 2082951896;
assign addr[27733]= 2100237377;
assign addr[27734]= 2114858546;
assign addr[27735]= 2126796855;
assign addr[27736]= 2136037160;
assign addr[27737]= 2142567738;
assign addr[27738]= 2146380306;
assign addr[27739]= 2147470025;
assign addr[27740]= 2145835515;
assign addr[27741]= 2141478848;
assign addr[27742]= 2134405552;
assign addr[27743]= 2124624598;
assign addr[27744]= 2112148396;
assign addr[27745]= 2096992772;
assign addr[27746]= 2079176953;
assign addr[27747]= 2058723538;
assign addr[27748]= 2035658475;
assign addr[27749]= 2010011024;
assign addr[27750]= 1981813720;
assign addr[27751]= 1951102334;
assign addr[27752]= 1917915825;
assign addr[27753]= 1882296293;
assign addr[27754]= 1844288924;
assign addr[27755]= 1803941934;
assign addr[27756]= 1761306505;
assign addr[27757]= 1716436725;
assign addr[27758]= 1669389513;
assign addr[27759]= 1620224553;
assign addr[27760]= 1569004214;
assign addr[27761]= 1515793473;
assign addr[27762]= 1460659832;
assign addr[27763]= 1403673233;
assign addr[27764]= 1344905966;
assign addr[27765]= 1284432584;
assign addr[27766]= 1222329801;
assign addr[27767]= 1158676398;
assign addr[27768]= 1093553126;
assign addr[27769]= 1027042599;
assign addr[27770]= 959229189;
assign addr[27771]= 890198924;
assign addr[27772]= 820039373;
assign addr[27773]= 748839539;
assign addr[27774]= 676689746;
assign addr[27775]= 603681519;
assign addr[27776]= 529907477;
assign addr[27777]= 455461206;
assign addr[27778]= 380437148;
assign addr[27779]= 304930476;
assign addr[27780]= 229036977;
assign addr[27781]= 152852926;
assign addr[27782]= 76474970;
assign addr[27783]= 0;
assign addr[27784]= -76474970;
assign addr[27785]= -152852926;
assign addr[27786]= -229036977;
assign addr[27787]= -304930476;
assign addr[27788]= -380437148;
assign addr[27789]= -455461206;
assign addr[27790]= -529907477;
assign addr[27791]= -603681519;
assign addr[27792]= -676689746;
assign addr[27793]= -748839539;
assign addr[27794]= -820039373;
assign addr[27795]= -890198924;
assign addr[27796]= -959229189;
assign addr[27797]= -1027042599;
assign addr[27798]= -1093553126;
assign addr[27799]= -1158676398;
assign addr[27800]= -1222329801;
assign addr[27801]= -1284432584;
assign addr[27802]= -1344905966;
assign addr[27803]= -1403673233;
assign addr[27804]= -1460659832;
assign addr[27805]= -1515793473;
assign addr[27806]= -1569004214;
assign addr[27807]= -1620224553;
assign addr[27808]= -1669389513;
assign addr[27809]= -1716436725;
assign addr[27810]= -1761306505;
assign addr[27811]= -1803941934;
assign addr[27812]= -1844288924;
assign addr[27813]= -1882296293;
assign addr[27814]= -1917915825;
assign addr[27815]= -1951102334;
assign addr[27816]= -1981813720;
assign addr[27817]= -2010011024;
assign addr[27818]= -2035658475;
assign addr[27819]= -2058723538;
assign addr[27820]= -2079176953;
assign addr[27821]= -2096992772;
assign addr[27822]= -2112148396;
assign addr[27823]= -2124624598;
assign addr[27824]= -2134405552;
assign addr[27825]= -2141478848;
assign addr[27826]= -2145835515;
assign addr[27827]= -2147470025;
assign addr[27828]= -2146380306;
assign addr[27829]= -2142567738;
assign addr[27830]= -2136037160;
assign addr[27831]= -2126796855;
assign addr[27832]= -2114858546;
assign addr[27833]= -2100237377;
assign addr[27834]= -2082951896;
assign addr[27835]= -2063024031;
assign addr[27836]= -2040479063;
assign addr[27837]= -2015345591;
assign addr[27838]= -1987655498;
assign addr[27839]= -1957443913;
assign addr[27840]= -1924749160;
assign addr[27841]= -1889612716;
assign addr[27842]= -1852079154;
assign addr[27843]= -1812196087;
assign addr[27844]= -1770014111;
assign addr[27845]= -1725586737;
assign addr[27846]= -1678970324;
assign addr[27847]= -1630224009;
assign addr[27848]= -1579409630;
assign addr[27849]= -1526591649;
assign addr[27850]= -1471837070;
assign addr[27851]= -1415215352;
assign addr[27852]= -1356798326;
assign addr[27853]= -1296660098;
assign addr[27854]= -1234876957;
assign addr[27855]= -1171527280;
assign addr[27856]= -1106691431;
assign addr[27857]= -1040451659;
assign addr[27858]= -972891995;
assign addr[27859]= -904098143;
assign addr[27860]= -834157373;
assign addr[27861]= -763158411;
assign addr[27862]= -691191324;
assign addr[27863]= -618347408;
assign addr[27864]= -544719071;
assign addr[27865]= -470399716;
assign addr[27866]= -395483624;
assign addr[27867]= -320065829;
assign addr[27868]= -244242007;
assign addr[27869]= -168108346;
assign addr[27870]= -91761426;
assign addr[27871]= -15298099;
assign addr[27872]= 61184634;
assign addr[27873]= 137589750;
assign addr[27874]= 213820322;
assign addr[27875]= 289779648;
assign addr[27876]= 365371365;
assign addr[27877]= 440499581;
assign addr[27878]= 515068990;
assign addr[27879]= 588984994;
assign addr[27880]= 662153826;
assign addr[27881]= 734482665;
assign addr[27882]= 805879757;
assign addr[27883]= 876254528;
assign addr[27884]= 945517704;
assign addr[27885]= 1013581418;
assign addr[27886]= 1080359326;
assign addr[27887]= 1145766716;
assign addr[27888]= 1209720613;
assign addr[27889]= 1272139887;
assign addr[27890]= 1332945355;
assign addr[27891]= 1392059879;
assign addr[27892]= 1449408469;
assign addr[27893]= 1504918373;
assign addr[27894]= 1558519173;
assign addr[27895]= 1610142873;
assign addr[27896]= 1659723983;
assign addr[27897]= 1707199606;
assign addr[27898]= 1752509516;
assign addr[27899]= 1795596234;
assign addr[27900]= 1836405100;
assign addr[27901]= 1874884346;
assign addr[27902]= 1910985158;
assign addr[27903]= 1944661739;
assign addr[27904]= 1975871368;
assign addr[27905]= 2004574453;
assign addr[27906]= 2030734582;
assign addr[27907]= 2054318569;
assign addr[27908]= 2075296495;
assign addr[27909]= 2093641749;
assign addr[27910]= 2109331059;
assign addr[27911]= 2122344521;
assign addr[27912]= 2132665626;
assign addr[27913]= 2140281282;
assign addr[27914]= 2145181827;
assign addr[27915]= 2147361045;
assign addr[27916]= 2146816171;
assign addr[27917]= 2143547897;
assign addr[27918]= 2137560369;
assign addr[27919]= 2128861181;
assign addr[27920]= 2117461370;
assign addr[27921]= 2103375398;
assign addr[27922]= 2086621133;
assign addr[27923]= 2067219829;
assign addr[27924]= 2045196100;
assign addr[27925]= 2020577882;
assign addr[27926]= 1993396407;
assign addr[27927]= 1963686155;
assign addr[27928]= 1931484818;
assign addr[27929]= 1896833245;
assign addr[27930]= 1859775393;
assign addr[27931]= 1820358275;
assign addr[27932]= 1778631892;
assign addr[27933]= 1734649179;
assign addr[27934]= 1688465931;
assign addr[27935]= 1640140734;
assign addr[27936]= 1589734894;
assign addr[27937]= 1537312353;
assign addr[27938]= 1482939614;
assign addr[27939]= 1426685652;
assign addr[27940]= 1368621831;
assign addr[27941]= 1308821808;
assign addr[27942]= 1247361445;
assign addr[27943]= 1184318708;
assign addr[27944]= 1119773573;
assign addr[27945]= 1053807919;
assign addr[27946]= 986505429;
assign addr[27947]= 917951481;
assign addr[27948]= 848233042;
assign addr[27949]= 777438554;
assign addr[27950]= 705657826;
assign addr[27951]= 632981917;
assign addr[27952]= 559503022;
assign addr[27953]= 485314355;
assign addr[27954]= 410510029;
assign addr[27955]= 335184940;
assign addr[27956]= 259434643;
assign addr[27957]= 183355234;
assign addr[27958]= 107043224;
assign addr[27959]= 30595422;
assign addr[27960]= -45891193;
assign addr[27961]= -122319591;
assign addr[27962]= -198592817;
assign addr[27963]= -274614114;
assign addr[27964]= -350287041;
assign addr[27965]= -425515602;
assign addr[27966]= -500204365;
assign addr[27967]= -574258580;
assign addr[27968]= -647584304;
assign addr[27969]= -720088517;
assign addr[27970]= -791679244;
assign addr[27971]= -862265664;
assign addr[27972]= -931758235;
assign addr[27973]= -1000068799;
assign addr[27974]= -1067110699;
assign addr[27975]= -1132798888;
assign addr[27976]= -1197050035;
assign addr[27977]= -1259782632;
assign addr[27978]= -1320917099;
assign addr[27979]= -1380375881;
assign addr[27980]= -1438083551;
assign addr[27981]= -1493966902;
assign addr[27982]= -1547955041;
assign addr[27983]= -1599979481;
assign addr[27984]= -1649974225;
assign addr[27985]= -1697875851;
assign addr[27986]= -1743623590;
assign addr[27987]= -1787159411;
assign addr[27988]= -1828428082;
assign addr[27989]= -1867377253;
assign addr[27990]= -1903957513;
assign addr[27991]= -1938122457;
assign addr[27992]= -1969828744;
assign addr[27993]= -1999036154;
assign addr[27994]= -2025707632;
assign addr[27995]= -2049809346;
assign addr[27996]= -2071310720;
assign addr[27997]= -2090184478;
assign addr[27998]= -2106406677;
assign addr[27999]= -2119956737;
assign addr[28000]= -2130817471;
assign addr[28001]= -2138975100;
assign addr[28002]= -2144419275;
assign addr[28003]= -2147143090;
assign addr[28004]= -2147143090;
assign addr[28005]= -2144419275;
assign addr[28006]= -2138975100;
assign addr[28007]= -2130817471;
assign addr[28008]= -2119956737;
assign addr[28009]= -2106406677;
assign addr[28010]= -2090184478;
assign addr[28011]= -2071310720;
assign addr[28012]= -2049809346;
assign addr[28013]= -2025707632;
assign addr[28014]= -1999036154;
assign addr[28015]= -1969828744;
assign addr[28016]= -1938122457;
assign addr[28017]= -1903957513;
assign addr[28018]= -1867377253;
assign addr[28019]= -1828428082;
assign addr[28020]= -1787159411;
assign addr[28021]= -1743623590;
assign addr[28022]= -1697875851;
assign addr[28023]= -1649974225;
assign addr[28024]= -1599979481;
assign addr[28025]= -1547955041;
assign addr[28026]= -1493966902;
assign addr[28027]= -1438083551;
assign addr[28028]= -1380375881;
assign addr[28029]= -1320917099;
assign addr[28030]= -1259782632;
assign addr[28031]= -1197050035;
assign addr[28032]= -1132798888;
assign addr[28033]= -1067110699;
assign addr[28034]= -1000068799;
assign addr[28035]= -931758235;
assign addr[28036]= -862265664;
assign addr[28037]= -791679244;
assign addr[28038]= -720088517;
assign addr[28039]= -647584304;
assign addr[28040]= -574258580;
assign addr[28041]= -500204365;
assign addr[28042]= -425515602;
assign addr[28043]= -350287041;
assign addr[28044]= -274614114;
assign addr[28045]= -198592817;
assign addr[28046]= -122319591;
assign addr[28047]= -45891193;
assign addr[28048]= 30595422;
assign addr[28049]= 107043224;
assign addr[28050]= 183355234;
assign addr[28051]= 259434643;
assign addr[28052]= 335184940;
assign addr[28053]= 410510029;
assign addr[28054]= 485314355;
assign addr[28055]= 559503022;
assign addr[28056]= 632981917;
assign addr[28057]= 705657826;
assign addr[28058]= 777438554;
assign addr[28059]= 848233042;
assign addr[28060]= 917951481;
assign addr[28061]= 986505429;
assign addr[28062]= 1053807919;
assign addr[28063]= 1119773573;
assign addr[28064]= 1184318708;
assign addr[28065]= 1247361445;
assign addr[28066]= 1308821808;
assign addr[28067]= 1368621831;
assign addr[28068]= 1426685652;
assign addr[28069]= 1482939614;
assign addr[28070]= 1537312353;
assign addr[28071]= 1589734894;
assign addr[28072]= 1640140734;
assign addr[28073]= 1688465931;
assign addr[28074]= 1734649179;
assign addr[28075]= 1778631892;
assign addr[28076]= 1820358275;
assign addr[28077]= 1859775393;
assign addr[28078]= 1896833245;
assign addr[28079]= 1931484818;
assign addr[28080]= 1963686155;
assign addr[28081]= 1993396407;
assign addr[28082]= 2020577882;
assign addr[28083]= 2045196100;
assign addr[28084]= 2067219829;
assign addr[28085]= 2086621133;
assign addr[28086]= 2103375398;
assign addr[28087]= 2117461370;
assign addr[28088]= 2128861181;
assign addr[28089]= 2137560369;
assign addr[28090]= 2143547897;
assign addr[28091]= 2146816171;
assign addr[28092]= 2147361045;
assign addr[28093]= 2145181827;
assign addr[28094]= 2140281282;
assign addr[28095]= 2132665626;
assign addr[28096]= 2122344521;
assign addr[28097]= 2109331059;
assign addr[28098]= 2093641749;
assign addr[28099]= 2075296495;
assign addr[28100]= 2054318569;
assign addr[28101]= 2030734582;
assign addr[28102]= 2004574453;
assign addr[28103]= 1975871368;
assign addr[28104]= 1944661739;
assign addr[28105]= 1910985158;
assign addr[28106]= 1874884346;
assign addr[28107]= 1836405100;
assign addr[28108]= 1795596234;
assign addr[28109]= 1752509516;
assign addr[28110]= 1707199606;
assign addr[28111]= 1659723983;
assign addr[28112]= 1610142873;
assign addr[28113]= 1558519173;
assign addr[28114]= 1504918373;
assign addr[28115]= 1449408469;
assign addr[28116]= 1392059879;
assign addr[28117]= 1332945355;
assign addr[28118]= 1272139887;
assign addr[28119]= 1209720613;
assign addr[28120]= 1145766716;
assign addr[28121]= 1080359326;
assign addr[28122]= 1013581418;
assign addr[28123]= 945517704;
assign addr[28124]= 876254528;
assign addr[28125]= 805879757;
assign addr[28126]= 734482665;
assign addr[28127]= 662153826;
assign addr[28128]= 588984994;
assign addr[28129]= 515068990;
assign addr[28130]= 440499581;
assign addr[28131]= 365371365;
assign addr[28132]= 289779648;
assign addr[28133]= 213820322;
assign addr[28134]= 137589750;
assign addr[28135]= 61184634;
assign addr[28136]= -15298099;
assign addr[28137]= -91761426;
assign addr[28138]= -168108346;
assign addr[28139]= -244242007;
assign addr[28140]= -320065829;
assign addr[28141]= -395483624;
assign addr[28142]= -470399716;
assign addr[28143]= -544719071;
assign addr[28144]= -618347408;
assign addr[28145]= -691191324;
assign addr[28146]= -763158411;
assign addr[28147]= -834157373;
assign addr[28148]= -904098143;
assign addr[28149]= -972891995;
assign addr[28150]= -1040451659;
assign addr[28151]= -1106691431;
assign addr[28152]= -1171527280;
assign addr[28153]= -1234876957;
assign addr[28154]= -1296660098;
assign addr[28155]= -1356798326;
assign addr[28156]= -1415215352;
assign addr[28157]= -1471837070;
assign addr[28158]= -1526591649;
assign addr[28159]= -1579409630;
assign addr[28160]= -1630224009;
assign addr[28161]= -1678970324;
assign addr[28162]= -1725586737;
assign addr[28163]= -1770014111;
assign addr[28164]= -1812196087;
assign addr[28165]= -1852079154;
assign addr[28166]= -1889612716;
assign addr[28167]= -1924749160;
assign addr[28168]= -1957443913;
assign addr[28169]= -1987655498;
assign addr[28170]= -2015345591;
assign addr[28171]= -2040479063;
assign addr[28172]= -2063024031;
assign addr[28173]= -2082951896;
assign addr[28174]= -2100237377;
assign addr[28175]= -2114858546;
assign addr[28176]= -2126796855;
assign addr[28177]= -2136037160;
assign addr[28178]= -2142567738;
assign addr[28179]= -2146380306;
assign addr[28180]= -2147470025;
assign addr[28181]= -2145835515;
assign addr[28182]= -2141478848;
assign addr[28183]= -2134405552;
assign addr[28184]= -2124624598;
assign addr[28185]= -2112148396;
assign addr[28186]= -2096992772;
assign addr[28187]= -2079176953;
assign addr[28188]= -2058723538;
assign addr[28189]= -2035658475;
assign addr[28190]= -2010011024;
assign addr[28191]= -1981813720;
assign addr[28192]= -1951102334;
assign addr[28193]= -1917915825;
assign addr[28194]= -1882296293;
assign addr[28195]= -1844288924;
assign addr[28196]= -1803941934;
assign addr[28197]= -1761306505;
assign addr[28198]= -1716436725;
assign addr[28199]= -1669389513;
assign addr[28200]= -1620224553;
assign addr[28201]= -1569004214;
assign addr[28202]= -1515793473;
assign addr[28203]= -1460659832;
assign addr[28204]= -1403673233;
assign addr[28205]= -1344905966;
assign addr[28206]= -1284432584;
assign addr[28207]= -1222329801;
assign addr[28208]= -1158676398;
assign addr[28209]= -1093553126;
assign addr[28210]= -1027042599;
assign addr[28211]= -959229189;
assign addr[28212]= -890198924;
assign addr[28213]= -820039373;
assign addr[28214]= -748839539;
assign addr[28215]= -676689746;
assign addr[28216]= -603681519;
assign addr[28217]= -529907477;
assign addr[28218]= -455461206;
assign addr[28219]= -380437148;
assign addr[28220]= -304930476;
assign addr[28221]= -229036977;
assign addr[28222]= -152852926;
assign addr[28223]= -76474970;
assign addr[28224]= 0;
assign addr[28225]= 76474970;
assign addr[28226]= 152852926;
assign addr[28227]= 229036977;
assign addr[28228]= 304930476;
assign addr[28229]= 380437148;
assign addr[28230]= 455461206;
assign addr[28231]= 529907477;
assign addr[28232]= 603681519;
assign addr[28233]= 676689746;
assign addr[28234]= 748839539;
assign addr[28235]= 820039373;
assign addr[28236]= 890198924;
assign addr[28237]= 959229189;
assign addr[28238]= 1027042599;
assign addr[28239]= 1093553126;
assign addr[28240]= 1158676398;
assign addr[28241]= 1222329801;
assign addr[28242]= 1284432584;
assign addr[28243]= 1344905966;
assign addr[28244]= 1403673233;
assign addr[28245]= 1460659832;
assign addr[28246]= 1515793473;
assign addr[28247]= 1569004214;
assign addr[28248]= 1620224553;
assign addr[28249]= 1669389513;
assign addr[28250]= 1716436725;
assign addr[28251]= 1761306505;
assign addr[28252]= 1803941934;
assign addr[28253]= 1844288924;
assign addr[28254]= 1882296293;
assign addr[28255]= 1917915825;
assign addr[28256]= 1951102334;
assign addr[28257]= 1981813720;
assign addr[28258]= 2010011024;
assign addr[28259]= 2035658475;
assign addr[28260]= 2058723538;
assign addr[28261]= 2079176953;
assign addr[28262]= 2096992772;
assign addr[28263]= 2112148396;
assign addr[28264]= 2124624598;
assign addr[28265]= 2134405552;
assign addr[28266]= 2141478848;
assign addr[28267]= 2145835515;
assign addr[28268]= 2147470025;
assign addr[28269]= 2146380306;
assign addr[28270]= 2142567738;
assign addr[28271]= 2136037160;
assign addr[28272]= 2126796855;
assign addr[28273]= 2114858546;
assign addr[28274]= 2100237377;
assign addr[28275]= 2082951896;
assign addr[28276]= 2063024031;
assign addr[28277]= 2040479063;
assign addr[28278]= 2015345591;
assign addr[28279]= 1987655498;
assign addr[28280]= 1957443913;
assign addr[28281]= 1924749160;
assign addr[28282]= 1889612716;
assign addr[28283]= 1852079154;
assign addr[28284]= 1812196087;
assign addr[28285]= 1770014111;
assign addr[28286]= 1725586737;
assign addr[28287]= 1678970324;
assign addr[28288]= 1630224009;
assign addr[28289]= 1579409630;
assign addr[28290]= 1526591649;
assign addr[28291]= 1471837070;
assign addr[28292]= 1415215352;
assign addr[28293]= 1356798326;
assign addr[28294]= 1296660098;
assign addr[28295]= 1234876957;
assign addr[28296]= 1171527280;
assign addr[28297]= 1106691431;
assign addr[28298]= 1040451659;
assign addr[28299]= 972891995;
assign addr[28300]= 904098143;
assign addr[28301]= 834157373;
assign addr[28302]= 763158411;
assign addr[28303]= 691191324;
assign addr[28304]= 618347408;
assign addr[28305]= 544719071;
assign addr[28306]= 470399716;
assign addr[28307]= 395483624;
assign addr[28308]= 320065829;
assign addr[28309]= 244242007;
assign addr[28310]= 168108346;
assign addr[28311]= 91761426;
assign addr[28312]= 15298099;
assign addr[28313]= -61184634;
assign addr[28314]= -137589750;
assign addr[28315]= -213820322;
assign addr[28316]= -289779648;
assign addr[28317]= -365371365;
assign addr[28318]= -440499581;
assign addr[28319]= -515068990;
assign addr[28320]= -588984994;
assign addr[28321]= -662153826;
assign addr[28322]= -734482665;
assign addr[28323]= -805879757;
assign addr[28324]= -876254528;
assign addr[28325]= -945517704;
assign addr[28326]= -1013581418;
assign addr[28327]= -1080359326;
assign addr[28328]= -1145766716;
assign addr[28329]= -1209720613;
assign addr[28330]= -1272139887;
assign addr[28331]= -1332945355;
assign addr[28332]= -1392059879;
assign addr[28333]= -1449408469;
assign addr[28334]= -1504918373;
assign addr[28335]= -1558519173;
assign addr[28336]= -1610142873;
assign addr[28337]= -1659723983;
assign addr[28338]= -1707199606;
assign addr[28339]= -1752509516;
assign addr[28340]= -1795596234;
assign addr[28341]= -1836405100;
assign addr[28342]= -1874884346;
assign addr[28343]= -1910985158;
assign addr[28344]= -1944661739;
assign addr[28345]= -1975871368;
assign addr[28346]= -2004574453;
assign addr[28347]= -2030734582;
assign addr[28348]= -2054318569;
assign addr[28349]= -2075296495;
assign addr[28350]= -2093641749;
assign addr[28351]= -2109331059;
assign addr[28352]= -2122344521;
assign addr[28353]= -2132665626;
assign addr[28354]= -2140281282;
assign addr[28355]= -2145181827;
assign addr[28356]= -2147361045;
assign addr[28357]= -2146816171;
assign addr[28358]= -2143547897;
assign addr[28359]= -2137560369;
assign addr[28360]= -2128861181;
assign addr[28361]= -2117461370;
assign addr[28362]= -2103375398;
assign addr[28363]= -2086621133;
assign addr[28364]= -2067219829;
assign addr[28365]= -2045196100;
assign addr[28366]= -2020577882;
assign addr[28367]= -1993396407;
assign addr[28368]= -1963686155;
assign addr[28369]= -1931484818;
assign addr[28370]= -1896833245;
assign addr[28371]= -1859775393;
assign addr[28372]= -1820358275;
assign addr[28373]= -1778631892;
assign addr[28374]= -1734649179;
assign addr[28375]= -1688465931;
assign addr[28376]= -1640140734;
assign addr[28377]= -1589734894;
assign addr[28378]= -1537312353;
assign addr[28379]= -1482939614;
assign addr[28380]= -1426685652;
assign addr[28381]= -1368621831;
assign addr[28382]= -1308821808;
assign addr[28383]= -1247361445;
assign addr[28384]= -1184318708;
assign addr[28385]= -1119773573;
assign addr[28386]= -1053807919;
assign addr[28387]= -986505429;
assign addr[28388]= -917951481;
assign addr[28389]= -848233042;
assign addr[28390]= -777438554;
assign addr[28391]= -705657826;
assign addr[28392]= -632981917;
assign addr[28393]= -559503022;
assign addr[28394]= -485314355;
assign addr[28395]= -410510029;
assign addr[28396]= -335184940;
assign addr[28397]= -259434643;
assign addr[28398]= -183355234;
assign addr[28399]= -107043224;
assign addr[28400]= -30595422;
assign addr[28401]= 45891193;
assign addr[28402]= 122319591;
assign addr[28403]= 198592817;
assign addr[28404]= 274614114;
assign addr[28405]= 350287041;
assign addr[28406]= 425515602;
assign addr[28407]= 500204365;
assign addr[28408]= 574258580;
assign addr[28409]= 647584304;
assign addr[28410]= 720088517;
assign addr[28411]= 791679244;
assign addr[28412]= 862265664;
assign addr[28413]= 931758235;
assign addr[28414]= 1000068799;
assign addr[28415]= 1067110699;
assign addr[28416]= 1132798888;
assign addr[28417]= 1197050035;
assign addr[28418]= 1259782632;
assign addr[28419]= 1320917099;
assign addr[28420]= 1380375881;
assign addr[28421]= 1438083551;
assign addr[28422]= 1493966902;
assign addr[28423]= 1547955041;
assign addr[28424]= 1599979481;
assign addr[28425]= 1649974225;
assign addr[28426]= 1697875851;
assign addr[28427]= 1743623590;
assign addr[28428]= 1787159411;
assign addr[28429]= 1828428082;
assign addr[28430]= 1867377253;
assign addr[28431]= 1903957513;
assign addr[28432]= 1938122457;
assign addr[28433]= 1969828744;
assign addr[28434]= 1999036154;
assign addr[28435]= 2025707632;
assign addr[28436]= 2049809346;
assign addr[28437]= 2071310720;
assign addr[28438]= 2090184478;
assign addr[28439]= 2106406677;
assign addr[28440]= 2119956737;
assign addr[28441]= 2130817471;
assign addr[28442]= 2138975100;
assign addr[28443]= 2144419275;
assign addr[28444]= 2147143090;
assign addr[28445]= 2147143090;
assign addr[28446]= 2144419275;
assign addr[28447]= 2138975100;
assign addr[28448]= 2130817471;
assign addr[28449]= 2119956737;
assign addr[28450]= 2106406677;
assign addr[28451]= 2090184478;
assign addr[28452]= 2071310720;
assign addr[28453]= 2049809346;
assign addr[28454]= 2025707632;
assign addr[28455]= 1999036154;
assign addr[28456]= 1969828744;
assign addr[28457]= 1938122457;
assign addr[28458]= 1903957513;
assign addr[28459]= 1867377253;
assign addr[28460]= 1828428082;
assign addr[28461]= 1787159411;
assign addr[28462]= 1743623590;
assign addr[28463]= 1697875851;
assign addr[28464]= 1649974225;
assign addr[28465]= 1599979481;
assign addr[28466]= 1547955041;
assign addr[28467]= 1493966902;
assign addr[28468]= 1438083551;
assign addr[28469]= 1380375881;
assign addr[28470]= 1320917099;
assign addr[28471]= 1259782632;
assign addr[28472]= 1197050035;
assign addr[28473]= 1132798888;
assign addr[28474]= 1067110699;
assign addr[28475]= 1000068799;
assign addr[28476]= 931758235;
assign addr[28477]= 862265664;
assign addr[28478]= 791679244;
assign addr[28479]= 720088517;
assign addr[28480]= 647584304;
assign addr[28481]= 574258580;
assign addr[28482]= 500204365;
assign addr[28483]= 425515602;
assign addr[28484]= 350287041;
assign addr[28485]= 274614114;
assign addr[28486]= 198592817;
assign addr[28487]= 122319591;
assign addr[28488]= 45891193;
assign addr[28489]= -30595422;
assign addr[28490]= -107043224;
assign addr[28491]= -183355234;
assign addr[28492]= -259434643;
assign addr[28493]= -335184940;
assign addr[28494]= -410510029;
assign addr[28495]= -485314355;
assign addr[28496]= -559503022;
assign addr[28497]= -632981917;
assign addr[28498]= -705657826;
assign addr[28499]= -777438554;
assign addr[28500]= -848233042;
assign addr[28501]= -917951481;
assign addr[28502]= -986505429;
assign addr[28503]= -1053807919;
assign addr[28504]= -1119773573;
assign addr[28505]= -1184318708;
assign addr[28506]= -1247361445;
assign addr[28507]= -1308821808;
assign addr[28508]= -1368621831;
assign addr[28509]= -1426685652;
assign addr[28510]= -1482939614;
assign addr[28511]= -1537312353;
assign addr[28512]= -1589734894;
assign addr[28513]= -1640140734;
assign addr[28514]= -1688465931;
assign addr[28515]= -1734649179;
assign addr[28516]= -1778631892;
assign addr[28517]= -1820358275;
assign addr[28518]= -1859775393;
assign addr[28519]= -1896833245;
assign addr[28520]= -1931484818;
assign addr[28521]= -1963686155;
assign addr[28522]= -1993396407;
assign addr[28523]= -2020577882;
assign addr[28524]= -2045196100;
assign addr[28525]= -2067219829;
assign addr[28526]= -2086621133;
assign addr[28527]= -2103375398;
assign addr[28528]= -2117461370;
assign addr[28529]= -2128861181;
assign addr[28530]= -2137560369;
assign addr[28531]= -2143547897;
assign addr[28532]= -2146816171;
assign addr[28533]= -2147361045;
assign addr[28534]= -2145181827;
assign addr[28535]= -2140281282;
assign addr[28536]= -2132665626;
assign addr[28537]= -2122344521;
assign addr[28538]= -2109331059;
assign addr[28539]= -2093641749;
assign addr[28540]= -2075296495;
assign addr[28541]= -2054318569;
assign addr[28542]= -2030734582;
assign addr[28543]= -2004574453;
assign addr[28544]= -1975871368;
assign addr[28545]= -1944661739;
assign addr[28546]= -1910985158;
assign addr[28547]= -1874884346;
assign addr[28548]= -1836405100;
assign addr[28549]= -1795596234;
assign addr[28550]= -1752509516;
assign addr[28551]= -1707199606;
assign addr[28552]= -1659723983;
assign addr[28553]= -1610142873;
assign addr[28554]= -1558519173;
assign addr[28555]= -1504918373;
assign addr[28556]= -1449408469;
assign addr[28557]= -1392059879;
assign addr[28558]= -1332945355;
assign addr[28559]= -1272139887;
assign addr[28560]= -1209720613;
assign addr[28561]= -1145766716;
assign addr[28562]= -1080359326;
assign addr[28563]= -1013581418;
assign addr[28564]= -945517704;
assign addr[28565]= -876254528;
assign addr[28566]= -805879757;
assign addr[28567]= -734482665;
assign addr[28568]= -662153826;
assign addr[28569]= -588984994;
assign addr[28570]= -515068990;
assign addr[28571]= -440499581;
assign addr[28572]= -365371365;
assign addr[28573]= -289779648;
assign addr[28574]= -213820322;
assign addr[28575]= -137589750;
assign addr[28576]= -61184634;
assign addr[28577]= 15298099;
assign addr[28578]= 91761426;
assign addr[28579]= 168108346;
assign addr[28580]= 244242007;
assign addr[28581]= 320065829;
assign addr[28582]= 395483624;
assign addr[28583]= 470399716;
assign addr[28584]= 544719071;
assign addr[28585]= 618347408;
assign addr[28586]= 691191324;
assign addr[28587]= 763158411;
assign addr[28588]= 834157373;
assign addr[28589]= 904098143;
assign addr[28590]= 972891995;
assign addr[28591]= 1040451659;
assign addr[28592]= 1106691431;
assign addr[28593]= 1171527280;
assign addr[28594]= 1234876957;
assign addr[28595]= 1296660098;
assign addr[28596]= 1356798326;
assign addr[28597]= 1415215352;
assign addr[28598]= 1471837070;
assign addr[28599]= 1526591649;
assign addr[28600]= 1579409630;
assign addr[28601]= 1630224009;
assign addr[28602]= 1678970324;
assign addr[28603]= 1725586737;
assign addr[28604]= 1770014111;
assign addr[28605]= 1812196087;
assign addr[28606]= 1852079154;
assign addr[28607]= 1889612716;
assign addr[28608]= 1924749160;
assign addr[28609]= 1957443913;
assign addr[28610]= 1987655498;
assign addr[28611]= 2015345591;
assign addr[28612]= 2040479063;
assign addr[28613]= 2063024031;
assign addr[28614]= 2082951896;
assign addr[28615]= 2100237377;
assign addr[28616]= 2114858546;
assign addr[28617]= 2126796855;
assign addr[28618]= 2136037160;
assign addr[28619]= 2142567738;
assign addr[28620]= 2146380306;
assign addr[28621]= 2147470025;
assign addr[28622]= 2145835515;
assign addr[28623]= 2141478848;
assign addr[28624]= 2134405552;
assign addr[28625]= 2124624598;
assign addr[28626]= 2112148396;
assign addr[28627]= 2096992772;
assign addr[28628]= 2079176953;
assign addr[28629]= 2058723538;
assign addr[28630]= 2035658475;
assign addr[28631]= 2010011024;
assign addr[28632]= 1981813720;
assign addr[28633]= 1951102334;
assign addr[28634]= 1917915825;
assign addr[28635]= 1882296293;
assign addr[28636]= 1844288924;
assign addr[28637]= 1803941934;
assign addr[28638]= 1761306505;
assign addr[28639]= 1716436725;
assign addr[28640]= 1669389513;
assign addr[28641]= 1620224553;
assign addr[28642]= 1569004214;
assign addr[28643]= 1515793473;
assign addr[28644]= 1460659832;
assign addr[28645]= 1403673233;
assign addr[28646]= 1344905966;
assign addr[28647]= 1284432584;
assign addr[28648]= 1222329801;
assign addr[28649]= 1158676398;
assign addr[28650]= 1093553126;
assign addr[28651]= 1027042599;
assign addr[28652]= 959229189;
assign addr[28653]= 890198924;
assign addr[28654]= 820039373;
assign addr[28655]= 748839539;
assign addr[28656]= 676689746;
assign addr[28657]= 603681519;
assign addr[28658]= 529907477;
assign addr[28659]= 455461206;
assign addr[28660]= 380437148;
assign addr[28661]= 304930476;
assign addr[28662]= 229036977;
assign addr[28663]= 152852926;
assign addr[28664]= 76474970;
assign addr[28665]= 0;
assign addr[28666]= -76474970;
assign addr[28667]= -152852926;
assign addr[28668]= -229036977;
assign addr[28669]= -304930476;
assign addr[28670]= -380437148;
assign addr[28671]= -455461206;
assign addr[28672]= -529907477;
assign addr[28673]= -603681519;
assign addr[28674]= -676689746;
assign addr[28675]= -748839539;
assign addr[28676]= -820039373;
assign addr[28677]= -890198924;
assign addr[28678]= -959229189;
assign addr[28679]= -1027042599;
assign addr[28680]= -1093553126;
assign addr[28681]= -1158676398;
assign addr[28682]= -1222329801;
assign addr[28683]= -1284432584;
assign addr[28684]= -1344905966;
assign addr[28685]= -1403673233;
assign addr[28686]= -1460659832;
assign addr[28687]= -1515793473;
assign addr[28688]= -1569004214;
assign addr[28689]= -1620224553;
assign addr[28690]= -1669389513;
assign addr[28691]= -1716436725;
assign addr[28692]= -1761306505;
assign addr[28693]= -1803941934;
assign addr[28694]= -1844288924;
assign addr[28695]= -1882296293;
assign addr[28696]= -1917915825;
assign addr[28697]= -1951102334;
assign addr[28698]= -1981813720;
assign addr[28699]= -2010011024;
assign addr[28700]= -2035658475;
assign addr[28701]= -2058723538;
assign addr[28702]= -2079176953;
assign addr[28703]= -2096992772;
assign addr[28704]= -2112148396;
assign addr[28705]= -2124624598;
assign addr[28706]= -2134405552;
assign addr[28707]= -2141478848;
assign addr[28708]= -2145835515;
assign addr[28709]= -2147470025;
assign addr[28710]= -2146380306;
assign addr[28711]= -2142567738;
assign addr[28712]= -2136037160;
assign addr[28713]= -2126796855;
assign addr[28714]= -2114858546;
assign addr[28715]= -2100237377;
assign addr[28716]= -2082951896;
assign addr[28717]= -2063024031;
assign addr[28718]= -2040479063;
assign addr[28719]= -2015345591;
assign addr[28720]= -1987655498;
assign addr[28721]= -1957443913;
assign addr[28722]= -1924749160;
assign addr[28723]= -1889612716;
assign addr[28724]= -1852079154;
assign addr[28725]= -1812196087;
assign addr[28726]= -1770014111;
assign addr[28727]= -1725586737;
assign addr[28728]= -1678970324;
assign addr[28729]= -1630224009;
assign addr[28730]= -1579409630;
assign addr[28731]= -1526591649;
assign addr[28732]= -1471837070;
assign addr[28733]= -1415215352;
assign addr[28734]= -1356798326;
assign addr[28735]= -1296660098;
assign addr[28736]= -1234876957;
assign addr[28737]= -1171527280;
assign addr[28738]= -1106691431;
assign addr[28739]= -1040451659;
assign addr[28740]= -972891995;
assign addr[28741]= -904098143;
assign addr[28742]= -834157373;
assign addr[28743]= -763158411;
assign addr[28744]= -691191324;
assign addr[28745]= -618347408;
assign addr[28746]= -544719071;
assign addr[28747]= -470399716;
assign addr[28748]= -395483624;
assign addr[28749]= -320065829;
assign addr[28750]= -244242007;
assign addr[28751]= -168108346;
assign addr[28752]= -91761426;
assign addr[28753]= -15298099;
assign addr[28754]= 61184634;
assign addr[28755]= 137589750;
assign addr[28756]= 213820322;
assign addr[28757]= 289779648;
assign addr[28758]= 365371365;
assign addr[28759]= 440499581;
assign addr[28760]= 515068990;
assign addr[28761]= 588984994;
assign addr[28762]= 662153826;
assign addr[28763]= 734482665;
assign addr[28764]= 805879757;
assign addr[28765]= 876254528;
assign addr[28766]= 945517704;
assign addr[28767]= 1013581418;
assign addr[28768]= 1080359326;
assign addr[28769]= 1145766716;
assign addr[28770]= 1209720613;
assign addr[28771]= 1272139887;
assign addr[28772]= 1332945355;
assign addr[28773]= 1392059879;
assign addr[28774]= 1449408469;
assign addr[28775]= 1504918373;
assign addr[28776]= 1558519173;
assign addr[28777]= 1610142873;
assign addr[28778]= 1659723983;
assign addr[28779]= 1707199606;
assign addr[28780]= 1752509516;
assign addr[28781]= 1795596234;
assign addr[28782]= 1836405100;
assign addr[28783]= 1874884346;
assign addr[28784]= 1910985158;
assign addr[28785]= 1944661739;
assign addr[28786]= 1975871368;
assign addr[28787]= 2004574453;
assign addr[28788]= 2030734582;
assign addr[28789]= 2054318569;
assign addr[28790]= 2075296495;
assign addr[28791]= 2093641749;
assign addr[28792]= 2109331059;
assign addr[28793]= 2122344521;
assign addr[28794]= 2132665626;
assign addr[28795]= 2140281282;
assign addr[28796]= 2145181827;
assign addr[28797]= 2147361045;
assign addr[28798]= 2146816171;
assign addr[28799]= 2143547897;
assign addr[28800]= 2137560369;
assign addr[28801]= 2128861181;
assign addr[28802]= 2117461370;
assign addr[28803]= 2103375398;
assign addr[28804]= 2086621133;
assign addr[28805]= 2067219829;
assign addr[28806]= 2045196100;
assign addr[28807]= 2020577882;
assign addr[28808]= 1993396407;
assign addr[28809]= 1963686155;
assign addr[28810]= 1931484818;
assign addr[28811]= 1896833245;
assign addr[28812]= 1859775393;
assign addr[28813]= 1820358275;
assign addr[28814]= 1778631892;
assign addr[28815]= 1734649179;
assign addr[28816]= 1688465931;
assign addr[28817]= 1640140734;
assign addr[28818]= 1589734894;
assign addr[28819]= 1537312353;
assign addr[28820]= 1482939614;
assign addr[28821]= 1426685652;
assign addr[28822]= 1368621831;
assign addr[28823]= 1308821808;
assign addr[28824]= 1247361445;
assign addr[28825]= 1184318708;
assign addr[28826]= 1119773573;
assign addr[28827]= 1053807919;
assign addr[28828]= 986505429;
assign addr[28829]= 917951481;
assign addr[28830]= 848233042;
assign addr[28831]= 777438554;
assign addr[28832]= 705657826;
assign addr[28833]= 632981917;
assign addr[28834]= 559503022;
assign addr[28835]= 485314355;
assign addr[28836]= 410510029;
assign addr[28837]= 335184940;
assign addr[28838]= 259434643;
assign addr[28839]= 183355234;
assign addr[28840]= 107043224;
assign addr[28841]= 30595422;
assign addr[28842]= -45891193;
assign addr[28843]= -122319591;
assign addr[28844]= -198592817;
assign addr[28845]= -274614114;
assign addr[28846]= -350287041;
assign addr[28847]= -425515602;
assign addr[28848]= -500204365;
assign addr[28849]= -574258580;
assign addr[28850]= -647584304;
assign addr[28851]= -720088517;
assign addr[28852]= -791679244;
assign addr[28853]= -862265664;
assign addr[28854]= -931758235;
assign addr[28855]= -1000068799;
assign addr[28856]= -1067110699;
assign addr[28857]= -1132798888;
assign addr[28858]= -1197050035;
assign addr[28859]= -1259782632;
assign addr[28860]= -1320917099;
assign addr[28861]= -1380375881;
assign addr[28862]= -1438083551;
assign addr[28863]= -1493966902;
assign addr[28864]= -1547955041;
assign addr[28865]= -1599979481;
assign addr[28866]= -1649974225;
assign addr[28867]= -1697875851;
assign addr[28868]= -1743623590;
assign addr[28869]= -1787159411;
assign addr[28870]= -1828428082;
assign addr[28871]= -1867377253;
assign addr[28872]= -1903957513;
assign addr[28873]= -1938122457;
assign addr[28874]= -1969828744;
assign addr[28875]= -1999036154;
assign addr[28876]= -2025707632;
assign addr[28877]= -2049809346;
assign addr[28878]= -2071310720;
assign addr[28879]= -2090184478;
assign addr[28880]= -2106406677;
assign addr[28881]= -2119956737;
assign addr[28882]= -2130817471;
assign addr[28883]= -2138975100;
assign addr[28884]= -2144419275;
assign addr[28885]= -2147143090;
assign addr[28886]= -2147143090;
assign addr[28887]= -2144419275;
assign addr[28888]= -2138975100;
assign addr[28889]= -2130817471;
assign addr[28890]= -2119956737;
assign addr[28891]= -2106406677;
assign addr[28892]= -2090184478;
assign addr[28893]= -2071310720;
assign addr[28894]= -2049809346;
assign addr[28895]= -2025707632;
assign addr[28896]= -1999036154;
assign addr[28897]= -1969828744;
assign addr[28898]= -1938122457;
assign addr[28899]= -1903957513;
assign addr[28900]= -1867377253;
assign addr[28901]= -1828428082;
assign addr[28902]= -1787159411;
assign addr[28903]= -1743623590;
assign addr[28904]= -1697875851;
assign addr[28905]= -1649974225;
assign addr[28906]= -1599979481;
assign addr[28907]= -1547955041;
assign addr[28908]= -1493966902;
assign addr[28909]= -1438083551;
assign addr[28910]= -1380375881;
assign addr[28911]= -1320917099;
assign addr[28912]= -1259782632;
assign addr[28913]= -1197050035;
assign addr[28914]= -1132798888;
assign addr[28915]= -1067110699;
assign addr[28916]= -1000068799;
assign addr[28917]= -931758235;
assign addr[28918]= -862265664;
assign addr[28919]= -791679244;
assign addr[28920]= -720088517;
assign addr[28921]= -647584304;
assign addr[28922]= -574258580;
assign addr[28923]= -500204365;
assign addr[28924]= -425515602;
assign addr[28925]= -350287041;
assign addr[28926]= -274614114;
assign addr[28927]= -198592817;
assign addr[28928]= -122319591;
assign addr[28929]= -45891193;
assign addr[28930]= 30595422;
assign addr[28931]= 107043224;
assign addr[28932]= 183355234;
assign addr[28933]= 259434643;
assign addr[28934]= 335184940;
assign addr[28935]= 410510029;
assign addr[28936]= 485314355;
assign addr[28937]= 559503022;
assign addr[28938]= 632981917;
assign addr[28939]= 705657826;
assign addr[28940]= 777438554;
assign addr[28941]= 848233042;
assign addr[28942]= 917951481;
assign addr[28943]= 986505429;
assign addr[28944]= 1053807919;
assign addr[28945]= 1119773573;
assign addr[28946]= 1184318708;
assign addr[28947]= 1247361445;
assign addr[28948]= 1308821808;
assign addr[28949]= 1368621831;
assign addr[28950]= 1426685652;
assign addr[28951]= 1482939614;
assign addr[28952]= 1537312353;
assign addr[28953]= 1589734894;
assign addr[28954]= 1640140734;
assign addr[28955]= 1688465931;
assign addr[28956]= 1734649179;
assign addr[28957]= 1778631892;
assign addr[28958]= 1820358275;
assign addr[28959]= 1859775393;
assign addr[28960]= 1896833245;
assign addr[28961]= 1931484818;
assign addr[28962]= 1963686155;
assign addr[28963]= 1993396407;
assign addr[28964]= 2020577882;
assign addr[28965]= 2045196100;
assign addr[28966]= 2067219829;
assign addr[28967]= 2086621133;
assign addr[28968]= 2103375398;
assign addr[28969]= 2117461370;
assign addr[28970]= 2128861181;
assign addr[28971]= 2137560369;
assign addr[28972]= 2143547897;
assign addr[28973]= 2146816171;
assign addr[28974]= 2147361045;
assign addr[28975]= 2145181827;
assign addr[28976]= 2140281282;
assign addr[28977]= 2132665626;
assign addr[28978]= 2122344521;
assign addr[28979]= 2109331059;
assign addr[28980]= 2093641749;
assign addr[28981]= 2075296495;
assign addr[28982]= 2054318569;
assign addr[28983]= 2030734582;
assign addr[28984]= 2004574453;
assign addr[28985]= 1975871368;
assign addr[28986]= 1944661739;
assign addr[28987]= 1910985158;
assign addr[28988]= 1874884346;
assign addr[28989]= 1836405100;
assign addr[28990]= 1795596234;
assign addr[28991]= 1752509516;
assign addr[28992]= 1707199606;
assign addr[28993]= 1659723983;
assign addr[28994]= 1610142873;
assign addr[28995]= 1558519173;
assign addr[28996]= 1504918373;
assign addr[28997]= 1449408469;
assign addr[28998]= 1392059879;
assign addr[28999]= 1332945355;
assign addr[29000]= 1272139887;
assign addr[29001]= 1209720613;
assign addr[29002]= 1145766716;
assign addr[29003]= 1080359326;
assign addr[29004]= 1013581418;
assign addr[29005]= 945517704;
assign addr[29006]= 876254528;
assign addr[29007]= 805879757;
assign addr[29008]= 734482665;
assign addr[29009]= 662153826;
assign addr[29010]= 588984994;
assign addr[29011]= 515068990;
assign addr[29012]= 440499581;
assign addr[29013]= 365371365;
assign addr[29014]= 289779648;
assign addr[29015]= 213820322;
assign addr[29016]= 137589750;
assign addr[29017]= 61184634;
assign addr[29018]= -15298099;
assign addr[29019]= -91761426;
assign addr[29020]= -168108346;
assign addr[29021]= -244242007;
assign addr[29022]= -320065829;
assign addr[29023]= -395483624;
assign addr[29024]= -470399716;
assign addr[29025]= -544719071;
assign addr[29026]= -618347408;
assign addr[29027]= -691191324;
assign addr[29028]= -763158411;
assign addr[29029]= -834157373;
assign addr[29030]= -904098143;
assign addr[29031]= -972891995;
assign addr[29032]= -1040451659;
assign addr[29033]= -1106691431;
assign addr[29034]= -1171527280;
assign addr[29035]= -1234876957;
assign addr[29036]= -1296660098;
assign addr[29037]= -1356798326;
assign addr[29038]= -1415215352;
assign addr[29039]= -1471837070;
assign addr[29040]= -1526591649;
assign addr[29041]= -1579409630;
assign addr[29042]= -1630224009;
assign addr[29043]= -1678970324;
assign addr[29044]= -1725586737;
assign addr[29045]= -1770014111;
assign addr[29046]= -1812196087;
assign addr[29047]= -1852079154;
assign addr[29048]= -1889612716;
assign addr[29049]= -1924749160;
assign addr[29050]= -1957443913;
assign addr[29051]= -1987655498;
assign addr[29052]= -2015345591;
assign addr[29053]= -2040479063;
assign addr[29054]= -2063024031;
assign addr[29055]= -2082951896;
assign addr[29056]= -2100237377;
assign addr[29057]= -2114858546;
assign addr[29058]= -2126796855;
assign addr[29059]= -2136037160;
assign addr[29060]= -2142567738;
assign addr[29061]= -2146380306;
assign addr[29062]= -2147470025;
assign addr[29063]= -2145835515;
assign addr[29064]= -2141478848;
assign addr[29065]= -2134405552;
assign addr[29066]= -2124624598;
assign addr[29067]= -2112148396;
assign addr[29068]= -2096992772;
assign addr[29069]= -2079176953;
assign addr[29070]= -2058723538;
assign addr[29071]= -2035658475;
assign addr[29072]= -2010011024;
assign addr[29073]= -1981813720;
assign addr[29074]= -1951102334;
assign addr[29075]= -1917915825;
assign addr[29076]= -1882296293;
assign addr[29077]= -1844288924;
assign addr[29078]= -1803941934;
assign addr[29079]= -1761306505;
assign addr[29080]= -1716436725;
assign addr[29081]= -1669389513;
assign addr[29082]= -1620224553;
assign addr[29083]= -1569004214;
assign addr[29084]= -1515793473;
assign addr[29085]= -1460659832;
assign addr[29086]= -1403673233;
assign addr[29087]= -1344905966;
assign addr[29088]= -1284432584;
assign addr[29089]= -1222329801;
assign addr[29090]= -1158676398;
assign addr[29091]= -1093553126;
assign addr[29092]= -1027042599;
assign addr[29093]= -959229189;
assign addr[29094]= -890198924;
assign addr[29095]= -820039373;
assign addr[29096]= -748839539;
assign addr[29097]= -676689746;
assign addr[29098]= -603681519;
assign addr[29099]= -529907477;
assign addr[29100]= -455461206;
assign addr[29101]= -380437148;
assign addr[29102]= -304930476;
assign addr[29103]= -229036977;
assign addr[29104]= -152852926;
assign addr[29105]= -76474970;
assign addr[29106]= 0;
assign addr[29107]= 76474970;
assign addr[29108]= 152852926;
assign addr[29109]= 229036977;
assign addr[29110]= 304930476;
assign addr[29111]= 380437148;
assign addr[29112]= 455461206;
assign addr[29113]= 529907477;
assign addr[29114]= 603681519;
assign addr[29115]= 676689746;
assign addr[29116]= 748839539;
assign addr[29117]= 820039373;
assign addr[29118]= 890198924;
assign addr[29119]= 959229189;
assign addr[29120]= 1027042599;
assign addr[29121]= 1093553126;
assign addr[29122]= 1158676398;
assign addr[29123]= 1222329801;
assign addr[29124]= 1284432584;
assign addr[29125]= 1344905966;
assign addr[29126]= 1403673233;
assign addr[29127]= 1460659832;
assign addr[29128]= 1515793473;
assign addr[29129]= 1569004214;
assign addr[29130]= 1620224553;
assign addr[29131]= 1669389513;
assign addr[29132]= 1716436725;
assign addr[29133]= 1761306505;
assign addr[29134]= 1803941934;
assign addr[29135]= 1844288924;
assign addr[29136]= 1882296293;
assign addr[29137]= 1917915825;
assign addr[29138]= 1951102334;
assign addr[29139]= 1981813720;
assign addr[29140]= 2010011024;
assign addr[29141]= 2035658475;
assign addr[29142]= 2058723538;
assign addr[29143]= 2079176953;
assign addr[29144]= 2096992772;
assign addr[29145]= 2112148396;
assign addr[29146]= 2124624598;
assign addr[29147]= 2134405552;
assign addr[29148]= 2141478848;
assign addr[29149]= 2145835515;
assign addr[29150]= 2147470025;
assign addr[29151]= 2146380306;
assign addr[29152]= 2142567738;
assign addr[29153]= 2136037160;
assign addr[29154]= 2126796855;
assign addr[29155]= 2114858546;
assign addr[29156]= 2100237377;
assign addr[29157]= 2082951896;
assign addr[29158]= 2063024031;
assign addr[29159]= 2040479063;
assign addr[29160]= 2015345591;
assign addr[29161]= 1987655498;
assign addr[29162]= 1957443913;
assign addr[29163]= 1924749160;
assign addr[29164]= 1889612716;
assign addr[29165]= 1852079154;
assign addr[29166]= 1812196087;
assign addr[29167]= 1770014111;
assign addr[29168]= 1725586737;
assign addr[29169]= 1678970324;
assign addr[29170]= 1630224009;
assign addr[29171]= 1579409630;
assign addr[29172]= 1526591649;
assign addr[29173]= 1471837070;
assign addr[29174]= 1415215352;
assign addr[29175]= 1356798326;
assign addr[29176]= 1296660098;
assign addr[29177]= 1234876957;
assign addr[29178]= 1171527280;
assign addr[29179]= 1106691431;
assign addr[29180]= 1040451659;
assign addr[29181]= 972891995;
assign addr[29182]= 904098143;
assign addr[29183]= 834157373;
assign addr[29184]= 763158411;
assign addr[29185]= 691191324;
assign addr[29186]= 618347408;
assign addr[29187]= 544719071;
assign addr[29188]= 470399716;
assign addr[29189]= 395483624;
assign addr[29190]= 320065829;
assign addr[29191]= 244242007;
assign addr[29192]= 168108346;
assign addr[29193]= 91761426;
assign addr[29194]= 15298099;
assign addr[29195]= -61184634;
assign addr[29196]= -137589750;
assign addr[29197]= -213820322;
assign addr[29198]= -289779648;
assign addr[29199]= -365371365;
assign addr[29200]= -440499581;
assign addr[29201]= -515068990;
assign addr[29202]= -588984994;
assign addr[29203]= -662153826;
assign addr[29204]= -734482665;
assign addr[29205]= -805879757;
assign addr[29206]= -876254528;
assign addr[29207]= -945517704;
assign addr[29208]= -1013581418;
assign addr[29209]= -1080359326;
assign addr[29210]= -1145766716;
assign addr[29211]= -1209720613;
assign addr[29212]= -1272139887;
assign addr[29213]= -1332945355;
assign addr[29214]= -1392059879;
assign addr[29215]= -1449408469;
assign addr[29216]= -1504918373;
assign addr[29217]= -1558519173;
assign addr[29218]= -1610142873;
assign addr[29219]= -1659723983;
assign addr[29220]= -1707199606;
assign addr[29221]= -1752509516;
assign addr[29222]= -1795596234;
assign addr[29223]= -1836405100;
assign addr[29224]= -1874884346;
assign addr[29225]= -1910985158;
assign addr[29226]= -1944661739;
assign addr[29227]= -1975871368;
assign addr[29228]= -2004574453;
assign addr[29229]= -2030734582;
assign addr[29230]= -2054318569;
assign addr[29231]= -2075296495;
assign addr[29232]= -2093641749;
assign addr[29233]= -2109331059;
assign addr[29234]= -2122344521;
assign addr[29235]= -2132665626;
assign addr[29236]= -2140281282;
assign addr[29237]= -2145181827;
assign addr[29238]= -2147361045;
assign addr[29239]= -2146816171;
assign addr[29240]= -2143547897;
assign addr[29241]= -2137560369;
assign addr[29242]= -2128861181;
assign addr[29243]= -2117461370;
assign addr[29244]= -2103375398;
assign addr[29245]= -2086621133;
assign addr[29246]= -2067219829;
assign addr[29247]= -2045196100;
assign addr[29248]= -2020577882;
assign addr[29249]= -1993396407;
assign addr[29250]= -1963686155;
assign addr[29251]= -1931484818;
assign addr[29252]= -1896833245;
assign addr[29253]= -1859775393;
assign addr[29254]= -1820358275;
assign addr[29255]= -1778631892;
assign addr[29256]= -1734649179;
assign addr[29257]= -1688465931;
assign addr[29258]= -1640140734;
assign addr[29259]= -1589734894;
assign addr[29260]= -1537312353;
assign addr[29261]= -1482939614;
assign addr[29262]= -1426685652;
assign addr[29263]= -1368621831;
assign addr[29264]= -1308821808;
assign addr[29265]= -1247361445;
assign addr[29266]= -1184318708;
assign addr[29267]= -1119773573;
assign addr[29268]= -1053807919;
assign addr[29269]= -986505429;
assign addr[29270]= -917951481;
assign addr[29271]= -848233042;
assign addr[29272]= -777438554;
assign addr[29273]= -705657826;
assign addr[29274]= -632981917;
assign addr[29275]= -559503022;
assign addr[29276]= -485314355;
assign addr[29277]= -410510029;
assign addr[29278]= -335184940;
assign addr[29279]= -259434643;
assign addr[29280]= -183355234;
assign addr[29281]= -107043224;
assign addr[29282]= -30595422;
assign addr[29283]= 45891193;
assign addr[29284]= 122319591;
assign addr[29285]= 198592817;
assign addr[29286]= 274614114;
assign addr[29287]= 350287041;
assign addr[29288]= 425515602;
assign addr[29289]= 500204365;
assign addr[29290]= 574258580;
assign addr[29291]= 647584304;
assign addr[29292]= 720088517;
assign addr[29293]= 791679244;
assign addr[29294]= 862265664;
assign addr[29295]= 931758235;
assign addr[29296]= 1000068799;
assign addr[29297]= 1067110699;
assign addr[29298]= 1132798888;
assign addr[29299]= 1197050035;
assign addr[29300]= 1259782632;
assign addr[29301]= 1320917099;
assign addr[29302]= 1380375881;
assign addr[29303]= 1438083551;
assign addr[29304]= 1493966902;
assign addr[29305]= 1547955041;
assign addr[29306]= 1599979481;
assign addr[29307]= 1649974225;
assign addr[29308]= 1697875851;
assign addr[29309]= 1743623590;
assign addr[29310]= 1787159411;
assign addr[29311]= 1828428082;
assign addr[29312]= 1867377253;
assign addr[29313]= 1903957513;
assign addr[29314]= 1938122457;
assign addr[29315]= 1969828744;
assign addr[29316]= 1999036154;
assign addr[29317]= 2025707632;
assign addr[29318]= 2049809346;
assign addr[29319]= 2071310720;
assign addr[29320]= 2090184478;
assign addr[29321]= 2106406677;
assign addr[29322]= 2119956737;
assign addr[29323]= 2130817471;
assign addr[29324]= 2138975100;
assign addr[29325]= 2144419275;
assign addr[29326]= 2147143090;
assign addr[29327]= 2147143090;
assign addr[29328]= 2144419275;
assign addr[29329]= 2138975100;
assign addr[29330]= 2130817471;
assign addr[29331]= 2119956737;
assign addr[29332]= 2106406677;
assign addr[29333]= 2090184478;
assign addr[29334]= 2071310720;
assign addr[29335]= 2049809346;
assign addr[29336]= 2025707632;
assign addr[29337]= 1999036154;
assign addr[29338]= 1969828744;
assign addr[29339]= 1938122457;
assign addr[29340]= 1903957513;
assign addr[29341]= 1867377253;
assign addr[29342]= 1828428082;
assign addr[29343]= 1787159411;
assign addr[29344]= 1743623590;
assign addr[29345]= 1697875851;
assign addr[29346]= 1649974225;
assign addr[29347]= 1599979481;
assign addr[29348]= 1547955041;
assign addr[29349]= 1493966902;
assign addr[29350]= 1438083551;
assign addr[29351]= 1380375881;
assign addr[29352]= 1320917099;
assign addr[29353]= 1259782632;
assign addr[29354]= 1197050035;
assign addr[29355]= 1132798888;
assign addr[29356]= 1067110699;
assign addr[29357]= 1000068799;
assign addr[29358]= 931758235;
assign addr[29359]= 862265664;
assign addr[29360]= 791679244;
assign addr[29361]= 720088517;
assign addr[29362]= 647584304;
assign addr[29363]= 574258580;
assign addr[29364]= 500204365;
assign addr[29365]= 425515602;
assign addr[29366]= 350287041;
assign addr[29367]= 274614114;
assign addr[29368]= 198592817;
assign addr[29369]= 122319591;
assign addr[29370]= 45891193;
assign addr[29371]= -30595422;
assign addr[29372]= -107043224;
assign addr[29373]= -183355234;
assign addr[29374]= -259434643;
assign addr[29375]= -335184940;
assign addr[29376]= -410510029;
assign addr[29377]= -485314355;
assign addr[29378]= -559503022;
assign addr[29379]= -632981917;
assign addr[29380]= -705657826;
assign addr[29381]= -777438554;
assign addr[29382]= -848233042;
assign addr[29383]= -917951481;
assign addr[29384]= -986505429;
assign addr[29385]= -1053807919;
assign addr[29386]= -1119773573;
assign addr[29387]= -1184318708;
assign addr[29388]= -1247361445;
assign addr[29389]= -1308821808;
assign addr[29390]= -1368621831;
assign addr[29391]= -1426685652;
assign addr[29392]= -1482939614;
assign addr[29393]= -1537312353;
assign addr[29394]= -1589734894;
assign addr[29395]= -1640140734;
assign addr[29396]= -1688465931;
assign addr[29397]= -1734649179;
assign addr[29398]= -1778631892;
assign addr[29399]= -1820358275;
assign addr[29400]= -1859775393;
assign addr[29401]= -1896833245;
assign addr[29402]= -1931484818;
assign addr[29403]= -1963686155;
assign addr[29404]= -1993396407;
assign addr[29405]= -2020577882;
assign addr[29406]= -2045196100;
assign addr[29407]= -2067219829;
assign addr[29408]= -2086621133;
assign addr[29409]= -2103375398;
assign addr[29410]= -2117461370;
assign addr[29411]= -2128861181;
assign addr[29412]= -2137560369;
assign addr[29413]= -2143547897;
assign addr[29414]= -2146816171;
assign addr[29415]= -2147361045;
assign addr[29416]= -2145181827;
assign addr[29417]= -2140281282;
assign addr[29418]= -2132665626;
assign addr[29419]= -2122344521;
assign addr[29420]= -2109331059;
assign addr[29421]= -2093641749;
assign addr[29422]= -2075296495;
assign addr[29423]= -2054318569;
assign addr[29424]= -2030734582;
assign addr[29425]= -2004574453;
assign addr[29426]= -1975871368;
assign addr[29427]= -1944661739;
assign addr[29428]= -1910985158;
assign addr[29429]= -1874884346;
assign addr[29430]= -1836405100;
assign addr[29431]= -1795596234;
assign addr[29432]= -1752509516;
assign addr[29433]= -1707199606;
assign addr[29434]= -1659723983;
assign addr[29435]= -1610142873;
assign addr[29436]= -1558519173;
assign addr[29437]= -1504918373;
assign addr[29438]= -1449408469;
assign addr[29439]= -1392059879;
assign addr[29440]= -1332945355;
assign addr[29441]= -1272139887;
assign addr[29442]= -1209720613;
assign addr[29443]= -1145766716;
assign addr[29444]= -1080359326;
assign addr[29445]= -1013581418;
assign addr[29446]= -945517704;
assign addr[29447]= -876254528;
assign addr[29448]= -805879757;
assign addr[29449]= -734482665;
assign addr[29450]= -662153826;
assign addr[29451]= -588984994;
assign addr[29452]= -515068990;
assign addr[29453]= -440499581;
assign addr[29454]= -365371365;
assign addr[29455]= -289779648;
assign addr[29456]= -213820322;
assign addr[29457]= -137589750;
assign addr[29458]= -61184634;
assign addr[29459]= 15298099;
assign addr[29460]= 91761426;
assign addr[29461]= 168108346;
assign addr[29462]= 244242007;
assign addr[29463]= 320065829;
assign addr[29464]= 395483624;
assign addr[29465]= 470399716;
assign addr[29466]= 544719071;
assign addr[29467]= 618347408;
assign addr[29468]= 691191324;
assign addr[29469]= 763158411;
assign addr[29470]= 834157373;
assign addr[29471]= 904098143;
assign addr[29472]= 972891995;
assign addr[29473]= 1040451659;
assign addr[29474]= 1106691431;
assign addr[29475]= 1171527280;
assign addr[29476]= 1234876957;
assign addr[29477]= 1296660098;
assign addr[29478]= 1356798326;
assign addr[29479]= 1415215352;
assign addr[29480]= 1471837070;
assign addr[29481]= 1526591649;
assign addr[29482]= 1579409630;
assign addr[29483]= 1630224009;
assign addr[29484]= 1678970324;
assign addr[29485]= 1725586737;
assign addr[29486]= 1770014111;
assign addr[29487]= 1812196087;
assign addr[29488]= 1852079154;
assign addr[29489]= 1889612716;
assign addr[29490]= 1924749160;
assign addr[29491]= 1957443913;
assign addr[29492]= 1987655498;
assign addr[29493]= 2015345591;
assign addr[29494]= 2040479063;
assign addr[29495]= 2063024031;
assign addr[29496]= 2082951896;
assign addr[29497]= 2100237377;
assign addr[29498]= 2114858546;
assign addr[29499]= 2126796855;
assign addr[29500]= 2136037160;
assign addr[29501]= 2142567738;
assign addr[29502]= 2146380306;
assign addr[29503]= 2147470025;
assign addr[29504]= 2145835515;
assign addr[29505]= 2141478848;
assign addr[29506]= 2134405552;
assign addr[29507]= 2124624598;
assign addr[29508]= 2112148396;
assign addr[29509]= 2096992772;
assign addr[29510]= 2079176953;
assign addr[29511]= 2058723538;
assign addr[29512]= 2035658475;
assign addr[29513]= 2010011024;
assign addr[29514]= 1981813720;
assign addr[29515]= 1951102334;
assign addr[29516]= 1917915825;
assign addr[29517]= 1882296293;
assign addr[29518]= 1844288924;
assign addr[29519]= 1803941934;
assign addr[29520]= 1761306505;
assign addr[29521]= 1716436725;
assign addr[29522]= 1669389513;
assign addr[29523]= 1620224553;
assign addr[29524]= 1569004214;
assign addr[29525]= 1515793473;
assign addr[29526]= 1460659832;
assign addr[29527]= 1403673233;
assign addr[29528]= 1344905966;
assign addr[29529]= 1284432584;
assign addr[29530]= 1222329801;
assign addr[29531]= 1158676398;
assign addr[29532]= 1093553126;
assign addr[29533]= 1027042599;
assign addr[29534]= 959229189;
assign addr[29535]= 890198924;
assign addr[29536]= 820039373;
assign addr[29537]= 748839539;
assign addr[29538]= 676689746;
assign addr[29539]= 603681519;
assign addr[29540]= 529907477;
assign addr[29541]= 455461206;
assign addr[29542]= 380437148;
assign addr[29543]= 304930476;
assign addr[29544]= 229036977;
assign addr[29545]= 152852926;
assign addr[29546]= 76474970;
assign addr[29547]= 0;
assign addr[29548]= -76474970;
assign addr[29549]= -152852926;
assign addr[29550]= -229036977;
assign addr[29551]= -304930476;
assign addr[29552]= -380437148;
assign addr[29553]= -455461206;
assign addr[29554]= -529907477;
assign addr[29555]= -603681519;
assign addr[29556]= -676689746;
assign addr[29557]= -748839539;
assign addr[29558]= -820039373;
assign addr[29559]= -890198924;
assign addr[29560]= -959229189;
assign addr[29561]= -1027042599;
assign addr[29562]= -1093553126;
assign addr[29563]= -1158676398;
assign addr[29564]= -1222329801;
assign addr[29565]= -1284432584;
assign addr[29566]= -1344905966;
assign addr[29567]= -1403673233;
assign addr[29568]= -1460659832;
assign addr[29569]= -1515793473;
assign addr[29570]= -1569004214;
assign addr[29571]= -1620224553;
assign addr[29572]= -1669389513;
assign addr[29573]= -1716436725;
assign addr[29574]= -1761306505;
assign addr[29575]= -1803941934;
assign addr[29576]= -1844288924;
assign addr[29577]= -1882296293;
assign addr[29578]= -1917915825;
assign addr[29579]= -1951102334;
assign addr[29580]= -1981813720;
assign addr[29581]= -2010011024;
assign addr[29582]= -2035658475;
assign addr[29583]= -2058723538;
assign addr[29584]= -2079176953;
assign addr[29585]= -2096992772;
assign addr[29586]= -2112148396;
assign addr[29587]= -2124624598;
assign addr[29588]= -2134405552;
assign addr[29589]= -2141478848;
assign addr[29590]= -2145835515;
assign addr[29591]= -2147470025;
assign addr[29592]= -2146380306;
assign addr[29593]= -2142567738;
assign addr[29594]= -2136037160;
assign addr[29595]= -2126796855;
assign addr[29596]= -2114858546;
assign addr[29597]= -2100237377;
assign addr[29598]= -2082951896;
assign addr[29599]= -2063024031;
assign addr[29600]= -2040479063;
assign addr[29601]= -2015345591;
assign addr[29602]= -1987655498;
assign addr[29603]= -1957443913;
assign addr[29604]= -1924749160;
assign addr[29605]= -1889612716;
assign addr[29606]= -1852079154;
assign addr[29607]= -1812196087;
assign addr[29608]= -1770014111;
assign addr[29609]= -1725586737;
assign addr[29610]= -1678970324;
assign addr[29611]= -1630224009;
assign addr[29612]= -1579409630;
assign addr[29613]= -1526591649;
assign addr[29614]= -1471837070;
assign addr[29615]= -1415215352;
assign addr[29616]= -1356798326;
assign addr[29617]= -1296660098;
assign addr[29618]= -1234876957;
assign addr[29619]= -1171527280;
assign addr[29620]= -1106691431;
assign addr[29621]= -1040451659;
assign addr[29622]= -972891995;
assign addr[29623]= -904098143;
assign addr[29624]= -834157373;
assign addr[29625]= -763158411;
assign addr[29626]= -691191324;
assign addr[29627]= -618347408;
assign addr[29628]= -544719071;
assign addr[29629]= -470399716;
assign addr[29630]= -395483624;
assign addr[29631]= -320065829;
assign addr[29632]= -244242007;
assign addr[29633]= -168108346;
assign addr[29634]= -91761426;
assign addr[29635]= -15298099;
assign addr[29636]= 61184634;
assign addr[29637]= 137589750;
assign addr[29638]= 213820322;
assign addr[29639]= 289779648;
assign addr[29640]= 365371365;
assign addr[29641]= 440499581;
assign addr[29642]= 515068990;
assign addr[29643]= 588984994;
assign addr[29644]= 662153826;
assign addr[29645]= 734482665;
assign addr[29646]= 805879757;
assign addr[29647]= 876254528;
assign addr[29648]= 945517704;
assign addr[29649]= 1013581418;
assign addr[29650]= 1080359326;
assign addr[29651]= 1145766716;
assign addr[29652]= 1209720613;
assign addr[29653]= 1272139887;
assign addr[29654]= 1332945355;
assign addr[29655]= 1392059879;
assign addr[29656]= 1449408469;
assign addr[29657]= 1504918373;
assign addr[29658]= 1558519173;
assign addr[29659]= 1610142873;
assign addr[29660]= 1659723983;
assign addr[29661]= 1707199606;
assign addr[29662]= 1752509516;
assign addr[29663]= 1795596234;
assign addr[29664]= 1836405100;
assign addr[29665]= 1874884346;
assign addr[29666]= 1910985158;
assign addr[29667]= 1944661739;
assign addr[29668]= 1975871368;
assign addr[29669]= 2004574453;
assign addr[29670]= 2030734582;
assign addr[29671]= 2054318569;
assign addr[29672]= 2075296495;
assign addr[29673]= 2093641749;
assign addr[29674]= 2109331059;
assign addr[29675]= 2122344521;
assign addr[29676]= 2132665626;
assign addr[29677]= 2140281282;
assign addr[29678]= 2145181827;
assign addr[29679]= 2147361045;
assign addr[29680]= 2146816171;
assign addr[29681]= 2143547897;
assign addr[29682]= 2137560369;
assign addr[29683]= 2128861181;
assign addr[29684]= 2117461370;
assign addr[29685]= 2103375398;
assign addr[29686]= 2086621133;
assign addr[29687]= 2067219829;
assign addr[29688]= 2045196100;
assign addr[29689]= 2020577882;
assign addr[29690]= 1993396407;
assign addr[29691]= 1963686155;
assign addr[29692]= 1931484818;
assign addr[29693]= 1896833245;
assign addr[29694]= 1859775393;
assign addr[29695]= 1820358275;
assign addr[29696]= 1778631892;
assign addr[29697]= 1734649179;
assign addr[29698]= 1688465931;
assign addr[29699]= 1640140734;
assign addr[29700]= 1589734894;
assign addr[29701]= 1537312353;
assign addr[29702]= 1482939614;
assign addr[29703]= 1426685652;
assign addr[29704]= 1368621831;
assign addr[29705]= 1308821808;
assign addr[29706]= 1247361445;
assign addr[29707]= 1184318708;
assign addr[29708]= 1119773573;
assign addr[29709]= 1053807919;
assign addr[29710]= 986505429;
assign addr[29711]= 917951481;
assign addr[29712]= 848233042;
assign addr[29713]= 777438554;
assign addr[29714]= 705657826;
assign addr[29715]= 632981917;
assign addr[29716]= 559503022;
assign addr[29717]= 485314355;
assign addr[29718]= 410510029;
assign addr[29719]= 335184940;
assign addr[29720]= 259434643;
assign addr[29721]= 183355234;
assign addr[29722]= 107043224;
assign addr[29723]= 30595422;
assign addr[29724]= -45891193;
assign addr[29725]= -122319591;
assign addr[29726]= -198592817;
assign addr[29727]= -274614114;
assign addr[29728]= -350287041;
assign addr[29729]= -425515602;
assign addr[29730]= -500204365;
assign addr[29731]= -574258580;
assign addr[29732]= -647584304;
assign addr[29733]= -720088517;
assign addr[29734]= -791679244;
assign addr[29735]= -862265664;
assign addr[29736]= -931758235;
assign addr[29737]= -1000068799;
assign addr[29738]= -1067110699;
assign addr[29739]= -1132798888;
assign addr[29740]= -1197050035;
assign addr[29741]= -1259782632;
assign addr[29742]= -1320917099;
assign addr[29743]= -1380375881;
assign addr[29744]= -1438083551;
assign addr[29745]= -1493966902;
assign addr[29746]= -1547955041;
assign addr[29747]= -1599979481;
assign addr[29748]= -1649974225;
assign addr[29749]= -1697875851;
assign addr[29750]= -1743623590;
assign addr[29751]= -1787159411;
assign addr[29752]= -1828428082;
assign addr[29753]= -1867377253;
assign addr[29754]= -1903957513;
assign addr[29755]= -1938122457;
assign addr[29756]= -1969828744;
assign addr[29757]= -1999036154;
assign addr[29758]= -2025707632;
assign addr[29759]= -2049809346;
assign addr[29760]= -2071310720;
assign addr[29761]= -2090184478;
assign addr[29762]= -2106406677;
assign addr[29763]= -2119956737;
assign addr[29764]= -2130817471;
assign addr[29765]= -2138975100;
assign addr[29766]= -2144419275;
assign addr[29767]= -2147143090;
assign addr[29768]= -2147143090;
assign addr[29769]= -2144419275;
assign addr[29770]= -2138975100;
assign addr[29771]= -2130817471;
assign addr[29772]= -2119956737;
assign addr[29773]= -2106406677;
assign addr[29774]= -2090184478;
assign addr[29775]= -2071310720;
assign addr[29776]= -2049809346;
assign addr[29777]= -2025707632;
assign addr[29778]= -1999036154;
assign addr[29779]= -1969828744;
assign addr[29780]= -1938122457;
assign addr[29781]= -1903957513;
assign addr[29782]= -1867377253;
assign addr[29783]= -1828428082;
assign addr[29784]= -1787159411;
assign addr[29785]= -1743623590;
assign addr[29786]= -1697875851;
assign addr[29787]= -1649974225;
assign addr[29788]= -1599979481;
assign addr[29789]= -1547955041;
assign addr[29790]= -1493966902;
assign addr[29791]= -1438083551;
assign addr[29792]= -1380375881;
assign addr[29793]= -1320917099;
assign addr[29794]= -1259782632;
assign addr[29795]= -1197050035;
assign addr[29796]= -1132798888;
assign addr[29797]= -1067110699;
assign addr[29798]= -1000068799;
assign addr[29799]= -931758235;
assign addr[29800]= -862265664;
assign addr[29801]= -791679244;
assign addr[29802]= -720088517;
assign addr[29803]= -647584304;
assign addr[29804]= -574258580;
assign addr[29805]= -500204365;
assign addr[29806]= -425515602;
assign addr[29807]= -350287041;
assign addr[29808]= -274614114;
assign addr[29809]= -198592817;
assign addr[29810]= -122319591;
assign addr[29811]= -45891193;
assign addr[29812]= 30595422;
assign addr[29813]= 107043224;
assign addr[29814]= 183355234;
assign addr[29815]= 259434643;
assign addr[29816]= 335184940;
assign addr[29817]= 410510029;
assign addr[29818]= 485314355;
assign addr[29819]= 559503022;
assign addr[29820]= 632981917;
assign addr[29821]= 705657826;
assign addr[29822]= 777438554;
assign addr[29823]= 848233042;
assign addr[29824]= 917951481;
assign addr[29825]= 986505429;
assign addr[29826]= 1053807919;
assign addr[29827]= 1119773573;
assign addr[29828]= 1184318708;
assign addr[29829]= 1247361445;
assign addr[29830]= 1308821808;
assign addr[29831]= 1368621831;
assign addr[29832]= 1426685652;
assign addr[29833]= 1482939614;
assign addr[29834]= 1537312353;
assign addr[29835]= 1589734894;
assign addr[29836]= 1640140734;
assign addr[29837]= 1688465931;
assign addr[29838]= 1734649179;
assign addr[29839]= 1778631892;
assign addr[29840]= 1820358275;
assign addr[29841]= 1859775393;
assign addr[29842]= 1896833245;
assign addr[29843]= 1931484818;
assign addr[29844]= 1963686155;
assign addr[29845]= 1993396407;
assign addr[29846]= 2020577882;
assign addr[29847]= 2045196100;
assign addr[29848]= 2067219829;
assign addr[29849]= 2086621133;
assign addr[29850]= 2103375398;
assign addr[29851]= 2117461370;
assign addr[29852]= 2128861181;
assign addr[29853]= 2137560369;
assign addr[29854]= 2143547897;
assign addr[29855]= 2146816171;
assign addr[29856]= 2147361045;
assign addr[29857]= 2145181827;
assign addr[29858]= 2140281282;
assign addr[29859]= 2132665626;
assign addr[29860]= 2122344521;
assign addr[29861]= 2109331059;
assign addr[29862]= 2093641749;
assign addr[29863]= 2075296495;
assign addr[29864]= 2054318569;
assign addr[29865]= 2030734582;
assign addr[29866]= 2004574453;
assign addr[29867]= 1975871368;
assign addr[29868]= 1944661739;
assign addr[29869]= 1910985158;
assign addr[29870]= 1874884346;
assign addr[29871]= 1836405100;
assign addr[29872]= 1795596234;
assign addr[29873]= 1752509516;
assign addr[29874]= 1707199606;
assign addr[29875]= 1659723983;
assign addr[29876]= 1610142873;
assign addr[29877]= 1558519173;
assign addr[29878]= 1504918373;
assign addr[29879]= 1449408469;
assign addr[29880]= 1392059879;
assign addr[29881]= 1332945355;
assign addr[29882]= 1272139887;
assign addr[29883]= 1209720613;
assign addr[29884]= 1145766716;
assign addr[29885]= 1080359326;
assign addr[29886]= 1013581418;
assign addr[29887]= 945517704;
assign addr[29888]= 876254528;
assign addr[29889]= 805879757;
assign addr[29890]= 734482665;
assign addr[29891]= 662153826;
assign addr[29892]= 588984994;
assign addr[29893]= 515068990;
assign addr[29894]= 440499581;
assign addr[29895]= 365371365;
assign addr[29896]= 289779648;
assign addr[29897]= 213820322;
assign addr[29898]= 137589750;
assign addr[29899]= 61184634;
assign addr[29900]= -15298099;
assign addr[29901]= -91761426;
assign addr[29902]= -168108346;
assign addr[29903]= -244242007;
assign addr[29904]= -320065829;
assign addr[29905]= -395483624;
assign addr[29906]= -470399716;
assign addr[29907]= -544719071;
assign addr[29908]= -618347408;
assign addr[29909]= -691191324;
assign addr[29910]= -763158411;
assign addr[29911]= -834157373;
assign addr[29912]= -904098143;
assign addr[29913]= -972891995;
assign addr[29914]= -1040451659;
assign addr[29915]= -1106691431;
assign addr[29916]= -1171527280;
assign addr[29917]= -1234876957;
assign addr[29918]= -1296660098;
assign addr[29919]= -1356798326;
assign addr[29920]= -1415215352;
assign addr[29921]= -1471837070;
assign addr[29922]= -1526591649;
assign addr[29923]= -1579409630;
assign addr[29924]= -1630224009;
assign addr[29925]= -1678970324;
assign addr[29926]= -1725586737;
assign addr[29927]= -1770014111;
assign addr[29928]= -1812196087;
assign addr[29929]= -1852079154;
assign addr[29930]= -1889612716;
assign addr[29931]= -1924749160;
assign addr[29932]= -1957443913;
assign addr[29933]= -1987655498;
assign addr[29934]= -2015345591;
assign addr[29935]= -2040479063;
assign addr[29936]= -2063024031;
assign addr[29937]= -2082951896;
assign addr[29938]= -2100237377;
assign addr[29939]= -2114858546;
assign addr[29940]= -2126796855;
assign addr[29941]= -2136037160;
assign addr[29942]= -2142567738;
assign addr[29943]= -2146380306;
assign addr[29944]= -2147470025;
assign addr[29945]= -2145835515;
assign addr[29946]= -2141478848;
assign addr[29947]= -2134405552;
assign addr[29948]= -2124624598;
assign addr[29949]= -2112148396;
assign addr[29950]= -2096992772;
assign addr[29951]= -2079176953;
assign addr[29952]= -2058723538;
assign addr[29953]= -2035658475;
assign addr[29954]= -2010011024;
assign addr[29955]= -1981813720;
assign addr[29956]= -1951102334;
assign addr[29957]= -1917915825;
assign addr[29958]= -1882296293;
assign addr[29959]= -1844288924;
assign addr[29960]= -1803941934;
assign addr[29961]= -1761306505;
assign addr[29962]= -1716436725;
assign addr[29963]= -1669389513;
assign addr[29964]= -1620224553;
assign addr[29965]= -1569004214;
assign addr[29966]= -1515793473;
assign addr[29967]= -1460659832;
assign addr[29968]= -1403673233;
assign addr[29969]= -1344905966;
assign addr[29970]= -1284432584;
assign addr[29971]= -1222329801;
assign addr[29972]= -1158676398;
assign addr[29973]= -1093553126;
assign addr[29974]= -1027042599;
assign addr[29975]= -959229189;
assign addr[29976]= -890198924;
assign addr[29977]= -820039373;
assign addr[29978]= -748839539;
assign addr[29979]= -676689746;
assign addr[29980]= -603681519;
assign addr[29981]= -529907477;
assign addr[29982]= -455461206;
assign addr[29983]= -380437148;
assign addr[29984]= -304930476;
assign addr[29985]= -229036977;
assign addr[29986]= -152852926;
assign addr[29987]= -76474970;
assign addr[29988]= 0;
assign addr[29989]= 76474970;
assign addr[29990]= 152852926;
assign addr[29991]= 229036977;
assign addr[29992]= 304930476;
assign addr[29993]= 380437148;
assign addr[29994]= 455461206;
assign addr[29995]= 529907477;
assign addr[29996]= 603681519;
assign addr[29997]= 676689746;
assign addr[29998]= 748839539;
assign addr[29999]= 820039373;
assign addr[30000]= 890198924;
assign addr[30001]= 959229189;
assign addr[30002]= 1027042599;
assign addr[30003]= 1093553126;
assign addr[30004]= 1158676398;
assign addr[30005]= 1222329801;
assign addr[30006]= 1284432584;
assign addr[30007]= 1344905966;
assign addr[30008]= 1403673233;
assign addr[30009]= 1460659832;
assign addr[30010]= 1515793473;
assign addr[30011]= 1569004214;
assign addr[30012]= 1620224553;
assign addr[30013]= 1669389513;
assign addr[30014]= 1716436725;
assign addr[30015]= 1761306505;
assign addr[30016]= 1803941934;
assign addr[30017]= 1844288924;
assign addr[30018]= 1882296293;
assign addr[30019]= 1917915825;
assign addr[30020]= 1951102334;
assign addr[30021]= 1981813720;
assign addr[30022]= 2010011024;
assign addr[30023]= 2035658475;
assign addr[30024]= 2058723538;
assign addr[30025]= 2079176953;
assign addr[30026]= 2096992772;
assign addr[30027]= 2112148396;
assign addr[30028]= 2124624598;
assign addr[30029]= 2134405552;
assign addr[30030]= 2141478848;
assign addr[30031]= 2145835515;
assign addr[30032]= 2147470025;
assign addr[30033]= 2146380306;
assign addr[30034]= 2142567738;
assign addr[30035]= 2136037160;
assign addr[30036]= 2126796855;
assign addr[30037]= 2114858546;
assign addr[30038]= 2100237377;
assign addr[30039]= 2082951896;
assign addr[30040]= 2063024031;
assign addr[30041]= 2040479063;
assign addr[30042]= 2015345591;
assign addr[30043]= 1987655498;
assign addr[30044]= 1957443913;
assign addr[30045]= 1924749160;
assign addr[30046]= 1889612716;
assign addr[30047]= 1852079154;
assign addr[30048]= 1812196087;
assign addr[30049]= 1770014111;
assign addr[30050]= 1725586737;
assign addr[30051]= 1678970324;
assign addr[30052]= 1630224009;
assign addr[30053]= 1579409630;
assign addr[30054]= 1526591649;
assign addr[30055]= 1471837070;
assign addr[30056]= 1415215352;
assign addr[30057]= 1356798326;
assign addr[30058]= 1296660098;
assign addr[30059]= 1234876957;
assign addr[30060]= 1171527280;
assign addr[30061]= 1106691431;
assign addr[30062]= 1040451659;
assign addr[30063]= 972891995;
assign addr[30064]= 904098143;
assign addr[30065]= 834157373;
assign addr[30066]= 763158411;
assign addr[30067]= 691191324;
assign addr[30068]= 618347408;
assign addr[30069]= 544719071;
assign addr[30070]= 470399716;
assign addr[30071]= 395483624;
assign addr[30072]= 320065829;
assign addr[30073]= 244242007;
assign addr[30074]= 168108346;
assign addr[30075]= 91761426;
assign addr[30076]= 15298099;
assign addr[30077]= -61184634;
assign addr[30078]= -137589750;
assign addr[30079]= -213820322;
assign addr[30080]= -289779648;
assign addr[30081]= -365371365;
assign addr[30082]= -440499581;
assign addr[30083]= -515068990;
assign addr[30084]= -588984994;
assign addr[30085]= -662153826;
assign addr[30086]= -734482665;
assign addr[30087]= -805879757;
assign addr[30088]= -876254528;
assign addr[30089]= -945517704;
assign addr[30090]= -1013581418;
assign addr[30091]= -1080359326;
assign addr[30092]= -1145766716;
assign addr[30093]= -1209720613;
assign addr[30094]= -1272139887;
assign addr[30095]= -1332945355;
assign addr[30096]= -1392059879;
assign addr[30097]= -1449408469;
assign addr[30098]= -1504918373;
assign addr[30099]= -1558519173;
assign addr[30100]= -1610142873;
assign addr[30101]= -1659723983;
assign addr[30102]= -1707199606;
assign addr[30103]= -1752509516;
assign addr[30104]= -1795596234;
assign addr[30105]= -1836405100;
assign addr[30106]= -1874884346;
assign addr[30107]= -1910985158;
assign addr[30108]= -1944661739;
assign addr[30109]= -1975871368;
assign addr[30110]= -2004574453;
assign addr[30111]= -2030734582;
assign addr[30112]= -2054318569;
assign addr[30113]= -2075296495;
assign addr[30114]= -2093641749;
assign addr[30115]= -2109331059;
assign addr[30116]= -2122344521;
assign addr[30117]= -2132665626;
assign addr[30118]= -2140281282;
assign addr[30119]= -2145181827;
assign addr[30120]= -2147361045;
assign addr[30121]= -2146816171;
assign addr[30122]= -2143547897;
assign addr[30123]= -2137560369;
assign addr[30124]= -2128861181;
assign addr[30125]= -2117461370;
assign addr[30126]= -2103375398;
assign addr[30127]= -2086621133;
assign addr[30128]= -2067219829;
assign addr[30129]= -2045196100;
assign addr[30130]= -2020577882;
assign addr[30131]= -1993396407;
assign addr[30132]= -1963686155;
assign addr[30133]= -1931484818;
assign addr[30134]= -1896833245;
assign addr[30135]= -1859775393;
assign addr[30136]= -1820358275;
assign addr[30137]= -1778631892;
assign addr[30138]= -1734649179;
assign addr[30139]= -1688465931;
assign addr[30140]= -1640140734;
assign addr[30141]= -1589734894;
assign addr[30142]= -1537312353;
assign addr[30143]= -1482939614;
assign addr[30144]= -1426685652;
assign addr[30145]= -1368621831;
assign addr[30146]= -1308821808;
assign addr[30147]= -1247361445;
assign addr[30148]= -1184318708;
assign addr[30149]= -1119773573;
assign addr[30150]= -1053807919;
assign addr[30151]= -986505429;
assign addr[30152]= -917951481;
assign addr[30153]= -848233042;
assign addr[30154]= -777438554;
assign addr[30155]= -705657826;
assign addr[30156]= -632981917;
assign addr[30157]= -559503022;
assign addr[30158]= -485314355;
assign addr[30159]= -410510029;
assign addr[30160]= -335184940;
assign addr[30161]= -259434643;
assign addr[30162]= -183355234;
assign addr[30163]= -107043224;
assign addr[30164]= -30595422;
assign addr[30165]= 45891193;
assign addr[30166]= 122319591;
assign addr[30167]= 198592817;
assign addr[30168]= 274614114;
assign addr[30169]= 350287041;
assign addr[30170]= 425515602;
assign addr[30171]= 500204365;
assign addr[30172]= 574258580;
assign addr[30173]= 647584304;
assign addr[30174]= 720088517;
assign addr[30175]= 791679244;
assign addr[30176]= 862265664;
assign addr[30177]= 931758235;
assign addr[30178]= 1000068799;
assign addr[30179]= 1067110699;
assign addr[30180]= 1132798888;
assign addr[30181]= 1197050035;
assign addr[30182]= 1259782632;
assign addr[30183]= 1320917099;
assign addr[30184]= 1380375881;
assign addr[30185]= 1438083551;
assign addr[30186]= 1493966902;
assign addr[30187]= 1547955041;
assign addr[30188]= 1599979481;
assign addr[30189]= 1649974225;
assign addr[30190]= 1697875851;
assign addr[30191]= 1743623590;
assign addr[30192]= 1787159411;
assign addr[30193]= 1828428082;
assign addr[30194]= 1867377253;
assign addr[30195]= 1903957513;
assign addr[30196]= 1938122457;
assign addr[30197]= 1969828744;
assign addr[30198]= 1999036154;
assign addr[30199]= 2025707632;
assign addr[30200]= 2049809346;
assign addr[30201]= 2071310720;
assign addr[30202]= 2090184478;
assign addr[30203]= 2106406677;
assign addr[30204]= 2119956737;
assign addr[30205]= 2130817471;
assign addr[30206]= 2138975100;
assign addr[30207]= 2144419275;
assign addr[30208]= 2147143090;
assign addr[30209]= 2147143090;
assign addr[30210]= 2144419275;
assign addr[30211]= 2138975100;
assign addr[30212]= 2130817471;
assign addr[30213]= 2119956737;
assign addr[30214]= 2106406677;
assign addr[30215]= 2090184478;
assign addr[30216]= 2071310720;
assign addr[30217]= 2049809346;
assign addr[30218]= 2025707632;
assign addr[30219]= 1999036154;
assign addr[30220]= 1969828744;
assign addr[30221]= 1938122457;
assign addr[30222]= 1903957513;
assign addr[30223]= 1867377253;
assign addr[30224]= 1828428082;
assign addr[30225]= 1787159411;
assign addr[30226]= 1743623590;
assign addr[30227]= 1697875851;
assign addr[30228]= 1649974225;
assign addr[30229]= 1599979481;
assign addr[30230]= 1547955041;
assign addr[30231]= 1493966902;
assign addr[30232]= 1438083551;
assign addr[30233]= 1380375881;
assign addr[30234]= 1320917099;
assign addr[30235]= 1259782632;
assign addr[30236]= 1197050035;
assign addr[30237]= 1132798888;
assign addr[30238]= 1067110699;
assign addr[30239]= 1000068799;
assign addr[30240]= 931758235;
assign addr[30241]= 862265664;
assign addr[30242]= 791679244;
assign addr[30243]= 720088517;
assign addr[30244]= 647584304;
assign addr[30245]= 574258580;
assign addr[30246]= 500204365;
assign addr[30247]= 425515602;
assign addr[30248]= 350287041;
assign addr[30249]= 274614114;
assign addr[30250]= 198592817;
assign addr[30251]= 122319591;
assign addr[30252]= 45891193;
assign addr[30253]= -30595422;
assign addr[30254]= -107043224;
assign addr[30255]= -183355234;
assign addr[30256]= -259434643;
assign addr[30257]= -335184940;
assign addr[30258]= -410510029;
assign addr[30259]= -485314355;
assign addr[30260]= -559503022;
assign addr[30261]= -632981917;
assign addr[30262]= -705657826;
assign addr[30263]= -777438554;
assign addr[30264]= -848233042;
assign addr[30265]= -917951481;
assign addr[30266]= -986505429;
assign addr[30267]= -1053807919;
assign addr[30268]= -1119773573;
assign addr[30269]= -1184318708;
assign addr[30270]= -1247361445;
assign addr[30271]= -1308821808;
assign addr[30272]= -1368621831;
assign addr[30273]= -1426685652;
assign addr[30274]= -1482939614;
assign addr[30275]= -1537312353;
assign addr[30276]= -1589734894;
assign addr[30277]= -1640140734;
assign addr[30278]= -1688465931;
assign addr[30279]= -1734649179;
assign addr[30280]= -1778631892;
assign addr[30281]= -1820358275;
assign addr[30282]= -1859775393;
assign addr[30283]= -1896833245;
assign addr[30284]= -1931484818;
assign addr[30285]= -1963686155;
assign addr[30286]= -1993396407;
assign addr[30287]= -2020577882;
assign addr[30288]= -2045196100;
assign addr[30289]= -2067219829;
assign addr[30290]= -2086621133;
assign addr[30291]= -2103375398;
assign addr[30292]= -2117461370;
assign addr[30293]= -2128861181;
assign addr[30294]= -2137560369;
assign addr[30295]= -2143547897;
assign addr[30296]= -2146816171;
assign addr[30297]= -2147361045;
assign addr[30298]= -2145181827;
assign addr[30299]= -2140281282;
assign addr[30300]= -2132665626;
assign addr[30301]= -2122344521;
assign addr[30302]= -2109331059;
assign addr[30303]= -2093641749;
assign addr[30304]= -2075296495;
assign addr[30305]= -2054318569;
assign addr[30306]= -2030734582;
assign addr[30307]= -2004574453;
assign addr[30308]= -1975871368;
assign addr[30309]= -1944661739;
assign addr[30310]= -1910985158;
assign addr[30311]= -1874884346;
assign addr[30312]= -1836405100;
assign addr[30313]= -1795596234;
assign addr[30314]= -1752509516;
assign addr[30315]= -1707199606;
assign addr[30316]= -1659723983;
assign addr[30317]= -1610142873;
assign addr[30318]= -1558519173;
assign addr[30319]= -1504918373;
assign addr[30320]= -1449408469;
assign addr[30321]= -1392059879;
assign addr[30322]= -1332945355;
assign addr[30323]= -1272139887;
assign addr[30324]= -1209720613;
assign addr[30325]= -1145766716;
assign addr[30326]= -1080359326;
assign addr[30327]= -1013581418;
assign addr[30328]= -945517704;
assign addr[30329]= -876254528;
assign addr[30330]= -805879757;
assign addr[30331]= -734482665;
assign addr[30332]= -662153826;
assign addr[30333]= -588984994;
assign addr[30334]= -515068990;
assign addr[30335]= -440499581;
assign addr[30336]= -365371365;
assign addr[30337]= -289779648;
assign addr[30338]= -213820322;
assign addr[30339]= -137589750;
assign addr[30340]= -61184634;
assign addr[30341]= 15298099;
assign addr[30342]= 91761426;
assign addr[30343]= 168108346;
assign addr[30344]= 244242007;
assign addr[30345]= 320065829;
assign addr[30346]= 395483624;
assign addr[30347]= 470399716;
assign addr[30348]= 544719071;
assign addr[30349]= 618347408;
assign addr[30350]= 691191324;
assign addr[30351]= 763158411;
assign addr[30352]= 834157373;
assign addr[30353]= 904098143;
assign addr[30354]= 972891995;
assign addr[30355]= 1040451659;
assign addr[30356]= 1106691431;
assign addr[30357]= 1171527280;
assign addr[30358]= 1234876957;
assign addr[30359]= 1296660098;
assign addr[30360]= 1356798326;
assign addr[30361]= 1415215352;
assign addr[30362]= 1471837070;
assign addr[30363]= 1526591649;
assign addr[30364]= 1579409630;
assign addr[30365]= 1630224009;
assign addr[30366]= 1678970324;
assign addr[30367]= 1725586737;
assign addr[30368]= 1770014111;
assign addr[30369]= 1812196087;
assign addr[30370]= 1852079154;
assign addr[30371]= 1889612716;
assign addr[30372]= 1924749160;
assign addr[30373]= 1957443913;
assign addr[30374]= 1987655498;
assign addr[30375]= 2015345591;
assign addr[30376]= 2040479063;
assign addr[30377]= 2063024031;
assign addr[30378]= 2082951896;
assign addr[30379]= 2100237377;
assign addr[30380]= 2114858546;
assign addr[30381]= 2126796855;
assign addr[30382]= 2136037160;
assign addr[30383]= 2142567738;
assign addr[30384]= 2146380306;
assign addr[30385]= 2147470025;
assign addr[30386]= 2145835515;
assign addr[30387]= 2141478848;
assign addr[30388]= 2134405552;
assign addr[30389]= 2124624598;
assign addr[30390]= 2112148396;
assign addr[30391]= 2096992772;
assign addr[30392]= 2079176953;
assign addr[30393]= 2058723538;
assign addr[30394]= 2035658475;
assign addr[30395]= 2010011024;
assign addr[30396]= 1981813720;
assign addr[30397]= 1951102334;
assign addr[30398]= 1917915825;
assign addr[30399]= 1882296293;
assign addr[30400]= 1844288924;
assign addr[30401]= 1803941934;
assign addr[30402]= 1761306505;
assign addr[30403]= 1716436725;
assign addr[30404]= 1669389513;
assign addr[30405]= 1620224553;
assign addr[30406]= 1569004214;
assign addr[30407]= 1515793473;
assign addr[30408]= 1460659832;
assign addr[30409]= 1403673233;
assign addr[30410]= 1344905966;
assign addr[30411]= 1284432584;
assign addr[30412]= 1222329801;
assign addr[30413]= 1158676398;
assign addr[30414]= 1093553126;
assign addr[30415]= 1027042599;
assign addr[30416]= 959229189;
assign addr[30417]= 890198924;
assign addr[30418]= 820039373;
assign addr[30419]= 748839539;
assign addr[30420]= 676689746;
assign addr[30421]= 603681519;
assign addr[30422]= 529907477;
assign addr[30423]= 455461206;
assign addr[30424]= 380437148;
assign addr[30425]= 304930476;
assign addr[30426]= 229036977;
assign addr[30427]= 152852926;
assign addr[30428]= 76474970;
assign addr[30429]= 0;
assign addr[30430]= -76474970;
assign addr[30431]= -152852926;
assign addr[30432]= -229036977;
assign addr[30433]= -304930476;
assign addr[30434]= -380437148;
assign addr[30435]= -455461206;
assign addr[30436]= -529907477;
assign addr[30437]= -603681519;
assign addr[30438]= -676689746;
assign addr[30439]= -748839539;
assign addr[30440]= -820039373;
assign addr[30441]= -890198924;
assign addr[30442]= -959229189;
assign addr[30443]= -1027042599;
assign addr[30444]= -1093553126;
assign addr[30445]= -1158676398;
assign addr[30446]= -1222329801;
assign addr[30447]= -1284432584;
assign addr[30448]= -1344905966;
assign addr[30449]= -1403673233;
assign addr[30450]= -1460659832;
assign addr[30451]= -1515793473;
assign addr[30452]= -1569004214;
assign addr[30453]= -1620224553;
assign addr[30454]= -1669389513;
assign addr[30455]= -1716436725;
assign addr[30456]= -1761306505;
assign addr[30457]= -1803941934;
assign addr[30458]= -1844288924;
assign addr[30459]= -1882296293;
assign addr[30460]= -1917915825;
assign addr[30461]= -1951102334;
assign addr[30462]= -1981813720;
assign addr[30463]= -2010011024;
assign addr[30464]= -2035658475;
assign addr[30465]= -2058723538;
assign addr[30466]= -2079176953;
assign addr[30467]= -2096992772;
assign addr[30468]= -2112148396;
assign addr[30469]= -2124624598;
assign addr[30470]= -2134405552;
assign addr[30471]= -2141478848;
assign addr[30472]= -2145835515;
assign addr[30473]= -2147470025;
assign addr[30474]= -2146380306;
assign addr[30475]= -2142567738;
assign addr[30476]= -2136037160;
assign addr[30477]= -2126796855;
assign addr[30478]= -2114858546;
assign addr[30479]= -2100237377;
assign addr[30480]= -2082951896;
assign addr[30481]= -2063024031;
assign addr[30482]= -2040479063;
assign addr[30483]= -2015345591;
assign addr[30484]= -1987655498;
assign addr[30485]= -1957443913;
assign addr[30486]= -1924749160;
assign addr[30487]= -1889612716;
assign addr[30488]= -1852079154;
assign addr[30489]= -1812196087;
assign addr[30490]= -1770014111;
assign addr[30491]= -1725586737;
assign addr[30492]= -1678970324;
assign addr[30493]= -1630224009;
assign addr[30494]= -1579409630;
assign addr[30495]= -1526591649;
assign addr[30496]= -1471837070;
assign addr[30497]= -1415215352;
assign addr[30498]= -1356798326;
assign addr[30499]= -1296660098;
assign addr[30500]= -1234876957;
assign addr[30501]= -1171527280;
assign addr[30502]= -1106691431;
assign addr[30503]= -1040451659;
assign addr[30504]= -972891995;
assign addr[30505]= -904098143;
assign addr[30506]= -834157373;
assign addr[30507]= -763158411;
assign addr[30508]= -691191324;
assign addr[30509]= -618347408;
assign addr[30510]= -544719071;
assign addr[30511]= -470399716;
assign addr[30512]= -395483624;
assign addr[30513]= -320065829;
assign addr[30514]= -244242007;
assign addr[30515]= -168108346;
assign addr[30516]= -91761426;
assign addr[30517]= -15298099;
assign addr[30518]= 61184634;
assign addr[30519]= 137589750;
assign addr[30520]= 213820322;
assign addr[30521]= 289779648;
assign addr[30522]= 365371365;
assign addr[30523]= 440499581;
assign addr[30524]= 515068990;
assign addr[30525]= 588984994;
assign addr[30526]= 662153826;
assign addr[30527]= 734482665;
assign addr[30528]= 805879757;
assign addr[30529]= 876254528;
assign addr[30530]= 945517704;
assign addr[30531]= 1013581418;
assign addr[30532]= 1080359326;
assign addr[30533]= 1145766716;
assign addr[30534]= 1209720613;
assign addr[30535]= 1272139887;
assign addr[30536]= 1332945355;
assign addr[30537]= 1392059879;
assign addr[30538]= 1449408469;
assign addr[30539]= 1504918373;
assign addr[30540]= 1558519173;
assign addr[30541]= 1610142873;
assign addr[30542]= 1659723983;
assign addr[30543]= 1707199606;
assign addr[30544]= 1752509516;
assign addr[30545]= 1795596234;
assign addr[30546]= 1836405100;
assign addr[30547]= 1874884346;
assign addr[30548]= 1910985158;
assign addr[30549]= 1944661739;
assign addr[30550]= 1975871368;
assign addr[30551]= 2004574453;
assign addr[30552]= 2030734582;
assign addr[30553]= 2054318569;
assign addr[30554]= 2075296495;
assign addr[30555]= 2093641749;
assign addr[30556]= 2109331059;
assign addr[30557]= 2122344521;
assign addr[30558]= 2132665626;
assign addr[30559]= 2140281282;
assign addr[30560]= 2145181827;
assign addr[30561]= 2147361045;
assign addr[30562]= 2146816171;
assign addr[30563]= 2143547897;
assign addr[30564]= 2137560369;
assign addr[30565]= 2128861181;
assign addr[30566]= 2117461370;
assign addr[30567]= 2103375398;
assign addr[30568]= 2086621133;
assign addr[30569]= 2067219829;
assign addr[30570]= 2045196100;
assign addr[30571]= 2020577882;
assign addr[30572]= 1993396407;
assign addr[30573]= 1963686155;
assign addr[30574]= 1931484818;
assign addr[30575]= 1896833245;
assign addr[30576]= 1859775393;
assign addr[30577]= 1820358275;
assign addr[30578]= 1778631892;
assign addr[30579]= 1734649179;
assign addr[30580]= 1688465931;
assign addr[30581]= 1640140734;
assign addr[30582]= 1589734894;
assign addr[30583]= 1537312353;
assign addr[30584]= 1482939614;
assign addr[30585]= 1426685652;
assign addr[30586]= 1368621831;
assign addr[30587]= 1308821808;
assign addr[30588]= 1247361445;
assign addr[30589]= 1184318708;
assign addr[30590]= 1119773573;
assign addr[30591]= 1053807919;
assign addr[30592]= 986505429;
assign addr[30593]= 917951481;
assign addr[30594]= 848233042;
assign addr[30595]= 777438554;
assign addr[30596]= 705657826;
assign addr[30597]= 632981917;
assign addr[30598]= 559503022;
assign addr[30599]= 485314355;
assign addr[30600]= 410510029;
assign addr[30601]= 335184940;
assign addr[30602]= 259434643;
assign addr[30603]= 183355234;
assign addr[30604]= 107043224;
assign addr[30605]= 30595422;
assign addr[30606]= -45891193;
assign addr[30607]= -122319591;
assign addr[30608]= -198592817;
assign addr[30609]= -274614114;
assign addr[30610]= -350287041;
assign addr[30611]= -425515602;
assign addr[30612]= -500204365;
assign addr[30613]= -574258580;
assign addr[30614]= -647584304;
assign addr[30615]= -720088517;
assign addr[30616]= -791679244;
assign addr[30617]= -862265664;
assign addr[30618]= -931758235;
assign addr[30619]= -1000068799;
assign addr[30620]= -1067110699;
assign addr[30621]= -1132798888;
assign addr[30622]= -1197050035;
assign addr[30623]= -1259782632;
assign addr[30624]= -1320917099;
assign addr[30625]= -1380375881;
assign addr[30626]= -1438083551;
assign addr[30627]= -1493966902;
assign addr[30628]= -1547955041;
assign addr[30629]= -1599979481;
assign addr[30630]= -1649974225;
assign addr[30631]= -1697875851;
assign addr[30632]= -1743623590;
assign addr[30633]= -1787159411;
assign addr[30634]= -1828428082;
assign addr[30635]= -1867377253;
assign addr[30636]= -1903957513;
assign addr[30637]= -1938122457;
assign addr[30638]= -1969828744;
assign addr[30639]= -1999036154;
assign addr[30640]= -2025707632;
assign addr[30641]= -2049809346;
assign addr[30642]= -2071310720;
assign addr[30643]= -2090184478;
assign addr[30644]= -2106406677;
assign addr[30645]= -2119956737;
assign addr[30646]= -2130817471;
assign addr[30647]= -2138975100;
assign addr[30648]= -2144419275;
assign addr[30649]= -2147143090;
assign addr[30650]= -2147143090;
assign addr[30651]= -2144419275;
assign addr[30652]= -2138975100;
assign addr[30653]= -2130817471;
assign addr[30654]= -2119956737;
assign addr[30655]= -2106406677;
assign addr[30656]= -2090184478;
assign addr[30657]= -2071310720;
assign addr[30658]= -2049809346;
assign addr[30659]= -2025707632;
assign addr[30660]= -1999036154;
assign addr[30661]= -1969828744;
assign addr[30662]= -1938122457;
assign addr[30663]= -1903957513;
assign addr[30664]= -1867377253;
assign addr[30665]= -1828428082;
assign addr[30666]= -1787159411;
assign addr[30667]= -1743623590;
assign addr[30668]= -1697875851;
assign addr[30669]= -1649974225;
assign addr[30670]= -1599979481;
assign addr[30671]= -1547955041;
assign addr[30672]= -1493966902;
assign addr[30673]= -1438083551;
assign addr[30674]= -1380375881;
assign addr[30675]= -1320917099;
assign addr[30676]= -1259782632;
assign addr[30677]= -1197050035;
assign addr[30678]= -1132798888;
assign addr[30679]= -1067110699;
assign addr[30680]= -1000068799;
assign addr[30681]= -931758235;
assign addr[30682]= -862265664;
assign addr[30683]= -791679244;
assign addr[30684]= -720088517;
assign addr[30685]= -647584304;
assign addr[30686]= -574258580;
assign addr[30687]= -500204365;
assign addr[30688]= -425515602;
assign addr[30689]= -350287041;
assign addr[30690]= -274614114;
assign addr[30691]= -198592817;
assign addr[30692]= -122319591;
assign addr[30693]= -45891193;
assign addr[30694]= 30595422;
assign addr[30695]= 107043224;
assign addr[30696]= 183355234;
assign addr[30697]= 259434643;
assign addr[30698]= 335184940;
assign addr[30699]= 410510029;
assign addr[30700]= 485314355;
assign addr[30701]= 559503022;
assign addr[30702]= 632981917;
assign addr[30703]= 705657826;
assign addr[30704]= 777438554;
assign addr[30705]= 848233042;
assign addr[30706]= 917951481;
assign addr[30707]= 986505429;
assign addr[30708]= 1053807919;
assign addr[30709]= 1119773573;
assign addr[30710]= 1184318708;
assign addr[30711]= 1247361445;
assign addr[30712]= 1308821808;
assign addr[30713]= 1368621831;
assign addr[30714]= 1426685652;
assign addr[30715]= 1482939614;
assign addr[30716]= 1537312353;
assign addr[30717]= 1589734894;
assign addr[30718]= 1640140734;
assign addr[30719]= 1688465931;
assign addr[30720]= 1734649179;
assign addr[30721]= 1778631892;
assign addr[30722]= 1820358275;
assign addr[30723]= 1859775393;
assign addr[30724]= 1896833245;
assign addr[30725]= 1931484818;
assign addr[30726]= 1963686155;
assign addr[30727]= 1993396407;
assign addr[30728]= 2020577882;
assign addr[30729]= 2045196100;
assign addr[30730]= 2067219829;
assign addr[30731]= 2086621133;
assign addr[30732]= 2103375398;
assign addr[30733]= 2117461370;
assign addr[30734]= 2128861181;
assign addr[30735]= 2137560369;
assign addr[30736]= 2143547897;
assign addr[30737]= 2146816171;
assign addr[30738]= 2147361045;
assign addr[30739]= 2145181827;
assign addr[30740]= 2140281282;
assign addr[30741]= 2132665626;
assign addr[30742]= 2122344521;
assign addr[30743]= 2109331059;
assign addr[30744]= 2093641749;
assign addr[30745]= 2075296495;
assign addr[30746]= 2054318569;
assign addr[30747]= 2030734582;
assign addr[30748]= 2004574453;
assign addr[30749]= 1975871368;
assign addr[30750]= 1944661739;
assign addr[30751]= 1910985158;
assign addr[30752]= 1874884346;
assign addr[30753]= 1836405100;
assign addr[30754]= 1795596234;
assign addr[30755]= 1752509516;
assign addr[30756]= 1707199606;
assign addr[30757]= 1659723983;
assign addr[30758]= 1610142873;
assign addr[30759]= 1558519173;
assign addr[30760]= 1504918373;
assign addr[30761]= 1449408469;
assign addr[30762]= 1392059879;
assign addr[30763]= 1332945355;
assign addr[30764]= 1272139887;
assign addr[30765]= 1209720613;
assign addr[30766]= 1145766716;
assign addr[30767]= 1080359326;
assign addr[30768]= 1013581418;
assign addr[30769]= 945517704;
assign addr[30770]= 876254528;
assign addr[30771]= 805879757;
assign addr[30772]= 734482665;
assign addr[30773]= 662153826;
assign addr[30774]= 588984994;
assign addr[30775]= 515068990;
assign addr[30776]= 440499581;
assign addr[30777]= 365371365;
assign addr[30778]= 289779648;
assign addr[30779]= 213820322;
assign addr[30780]= 137589750;
assign addr[30781]= 61184634;
assign addr[30782]= -15298099;
assign addr[30783]= -91761426;
assign addr[30784]= -168108346;
assign addr[30785]= -244242007;
assign addr[30786]= -320065829;
assign addr[30787]= -395483624;
assign addr[30788]= -470399716;
assign addr[30789]= -544719071;
assign addr[30790]= -618347408;
assign addr[30791]= -691191324;
assign addr[30792]= -763158411;
assign addr[30793]= -834157373;
assign addr[30794]= -904098143;
assign addr[30795]= -972891995;
assign addr[30796]= -1040451659;
assign addr[30797]= -1106691431;
assign addr[30798]= -1171527280;
assign addr[30799]= -1234876957;
assign addr[30800]= -1296660098;
assign addr[30801]= -1356798326;
assign addr[30802]= -1415215352;
assign addr[30803]= -1471837070;
assign addr[30804]= -1526591649;
assign addr[30805]= -1579409630;
assign addr[30806]= -1630224009;
assign addr[30807]= -1678970324;
assign addr[30808]= -1725586737;
assign addr[30809]= -1770014111;
assign addr[30810]= -1812196087;
assign addr[30811]= -1852079154;
assign addr[30812]= -1889612716;
assign addr[30813]= -1924749160;
assign addr[30814]= -1957443913;
assign addr[30815]= -1987655498;
assign addr[30816]= -2015345591;
assign addr[30817]= -2040479063;
assign addr[30818]= -2063024031;
assign addr[30819]= -2082951896;
assign addr[30820]= -2100237377;
assign addr[30821]= -2114858546;
assign addr[30822]= -2126796855;
assign addr[30823]= -2136037160;
assign addr[30824]= -2142567738;
assign addr[30825]= -2146380306;
assign addr[30826]= -2147470025;
assign addr[30827]= -2145835515;
assign addr[30828]= -2141478848;
assign addr[30829]= -2134405552;
assign addr[30830]= -2124624598;
assign addr[30831]= -2112148396;
assign addr[30832]= -2096992772;
assign addr[30833]= -2079176953;
assign addr[30834]= -2058723538;
assign addr[30835]= -2035658475;
assign addr[30836]= -2010011024;
assign addr[30837]= -1981813720;
assign addr[30838]= -1951102334;
assign addr[30839]= -1917915825;
assign addr[30840]= -1882296293;
assign addr[30841]= -1844288924;
assign addr[30842]= -1803941934;
assign addr[30843]= -1761306505;
assign addr[30844]= -1716436725;
assign addr[30845]= -1669389513;
assign addr[30846]= -1620224553;
assign addr[30847]= -1569004214;
assign addr[30848]= -1515793473;
assign addr[30849]= -1460659832;
assign addr[30850]= -1403673233;
assign addr[30851]= -1344905966;
assign addr[30852]= -1284432584;
assign addr[30853]= -1222329801;
assign addr[30854]= -1158676398;
assign addr[30855]= -1093553126;
assign addr[30856]= -1027042599;
assign addr[30857]= -959229189;
assign addr[30858]= -890198924;
assign addr[30859]= -820039373;
assign addr[30860]= -748839539;
assign addr[30861]= -676689746;
assign addr[30862]= -603681519;
assign addr[30863]= -529907477;
assign addr[30864]= -455461206;
assign addr[30865]= -380437148;
assign addr[30866]= -304930476;
assign addr[30867]= -229036977;
assign addr[30868]= -152852926;
assign addr[30869]= -76474970;
assign addr[30870]= 0;
assign addr[30871]= 76474970;
assign addr[30872]= 152852926;
assign addr[30873]= 229036977;
assign addr[30874]= 304930476;
assign addr[30875]= 380437148;
assign addr[30876]= 455461206;
assign addr[30877]= 529907477;
assign addr[30878]= 603681519;
assign addr[30879]= 676689746;
assign addr[30880]= 748839539;
assign addr[30881]= 820039373;
assign addr[30882]= 890198924;
assign addr[30883]= 959229189;
assign addr[30884]= 1027042599;
assign addr[30885]= 1093553126;
assign addr[30886]= 1158676398;
assign addr[30887]= 1222329801;
assign addr[30888]= 1284432584;
assign addr[30889]= 1344905966;
assign addr[30890]= 1403673233;
assign addr[30891]= 1460659832;
assign addr[30892]= 1515793473;
assign addr[30893]= 1569004214;
assign addr[30894]= 1620224553;
assign addr[30895]= 1669389513;
assign addr[30896]= 1716436725;
assign addr[30897]= 1761306505;
assign addr[30898]= 1803941934;
assign addr[30899]= 1844288924;
assign addr[30900]= 1882296293;
assign addr[30901]= 1917915825;
assign addr[30902]= 1951102334;
assign addr[30903]= 1981813720;
assign addr[30904]= 2010011024;
assign addr[30905]= 2035658475;
assign addr[30906]= 2058723538;
assign addr[30907]= 2079176953;
assign addr[30908]= 2096992772;
assign addr[30909]= 2112148396;
assign addr[30910]= 2124624598;
assign addr[30911]= 2134405552;
assign addr[30912]= 2141478848;
assign addr[30913]= 2145835515;
assign addr[30914]= 2147470025;
assign addr[30915]= 2146380306;
assign addr[30916]= 2142567738;
assign addr[30917]= 2136037160;
assign addr[30918]= 2126796855;
assign addr[30919]= 2114858546;
assign addr[30920]= 2100237377;
assign addr[30921]= 2082951896;
assign addr[30922]= 2063024031;
assign addr[30923]= 2040479063;
assign addr[30924]= 2015345591;
assign addr[30925]= 1987655498;
assign addr[30926]= 1957443913;
assign addr[30927]= 1924749160;
assign addr[30928]= 1889612716;
assign addr[30929]= 1852079154;
assign addr[30930]= 1812196087;
assign addr[30931]= 1770014111;
assign addr[30932]= 1725586737;
assign addr[30933]= 1678970324;
assign addr[30934]= 1630224009;
assign addr[30935]= 1579409630;
assign addr[30936]= 1526591649;
assign addr[30937]= 1471837070;
assign addr[30938]= 1415215352;
assign addr[30939]= 1356798326;
assign addr[30940]= 1296660098;
assign addr[30941]= 1234876957;
assign addr[30942]= 1171527280;
assign addr[30943]= 1106691431;
assign addr[30944]= 1040451659;
assign addr[30945]= 972891995;
assign addr[30946]= 904098143;
assign addr[30947]= 834157373;
assign addr[30948]= 763158411;
assign addr[30949]= 691191324;
assign addr[30950]= 618347408;
assign addr[30951]= 544719071;
assign addr[30952]= 470399716;
assign addr[30953]= 395483624;
assign addr[30954]= 320065829;
assign addr[30955]= 244242007;
assign addr[30956]= 168108346;
assign addr[30957]= 91761426;
assign addr[30958]= 15298099;
assign addr[30959]= -61184634;
assign addr[30960]= -137589750;
assign addr[30961]= -213820322;
assign addr[30962]= -289779648;
assign addr[30963]= -365371365;
assign addr[30964]= -440499581;
assign addr[30965]= -515068990;
assign addr[30966]= -588984994;
assign addr[30967]= -662153826;
assign addr[30968]= -734482665;
assign addr[30969]= -805879757;
assign addr[30970]= -876254528;
assign addr[30971]= -945517704;
assign addr[30972]= -1013581418;
assign addr[30973]= -1080359326;
assign addr[30974]= -1145766716;
assign addr[30975]= -1209720613;
assign addr[30976]= -1272139887;
assign addr[30977]= -1332945355;
assign addr[30978]= -1392059879;
assign addr[30979]= -1449408469;
assign addr[30980]= -1504918373;
assign addr[30981]= -1558519173;
assign addr[30982]= -1610142873;
assign addr[30983]= -1659723983;
assign addr[30984]= -1707199606;
assign addr[30985]= -1752509516;
assign addr[30986]= -1795596234;
assign addr[30987]= -1836405100;
assign addr[30988]= -1874884346;
assign addr[30989]= -1910985158;
assign addr[30990]= -1944661739;
assign addr[30991]= -1975871368;
assign addr[30992]= -2004574453;
assign addr[30993]= -2030734582;
assign addr[30994]= -2054318569;
assign addr[30995]= -2075296495;
assign addr[30996]= -2093641749;
assign addr[30997]= -2109331059;
assign addr[30998]= -2122344521;
assign addr[30999]= -2132665626;
assign addr[31000]= -2140281282;
assign addr[31001]= -2145181827;
assign addr[31002]= -2147361045;
assign addr[31003]= -2146816171;
assign addr[31004]= -2143547897;
assign addr[31005]= -2137560369;
assign addr[31006]= -2128861181;
assign addr[31007]= -2117461370;
assign addr[31008]= -2103375398;
assign addr[31009]= -2086621133;
assign addr[31010]= -2067219829;
assign addr[31011]= -2045196100;
assign addr[31012]= -2020577882;
assign addr[31013]= -1993396407;
assign addr[31014]= -1963686155;
assign addr[31015]= -1931484818;
assign addr[31016]= -1896833245;
assign addr[31017]= -1859775393;
assign addr[31018]= -1820358275;
assign addr[31019]= -1778631892;
assign addr[31020]= -1734649179;
assign addr[31021]= -1688465931;
assign addr[31022]= -1640140734;
assign addr[31023]= -1589734894;
assign addr[31024]= -1537312353;
assign addr[31025]= -1482939614;
assign addr[31026]= -1426685652;
assign addr[31027]= -1368621831;
assign addr[31028]= -1308821808;
assign addr[31029]= -1247361445;
assign addr[31030]= -1184318708;
assign addr[31031]= -1119773573;
assign addr[31032]= -1053807919;
assign addr[31033]= -986505429;
assign addr[31034]= -917951481;
assign addr[31035]= -848233042;
assign addr[31036]= -777438554;
assign addr[31037]= -705657826;
assign addr[31038]= -632981917;
assign addr[31039]= -559503022;
assign addr[31040]= -485314355;
assign addr[31041]= -410510029;
assign addr[31042]= -335184940;
assign addr[31043]= -259434643;
assign addr[31044]= -183355234;
assign addr[31045]= -107043224;
assign addr[31046]= -30595422;
assign addr[31047]= 45891193;
assign addr[31048]= 122319591;
assign addr[31049]= 198592817;
assign addr[31050]= 274614114;
assign addr[31051]= 350287041;
assign addr[31052]= 425515602;
assign addr[31053]= 500204365;
assign addr[31054]= 574258580;
assign addr[31055]= 647584304;
assign addr[31056]= 720088517;
assign addr[31057]= 791679244;
assign addr[31058]= 862265664;
assign addr[31059]= 931758235;
assign addr[31060]= 1000068799;
assign addr[31061]= 1067110699;
assign addr[31062]= 1132798888;
assign addr[31063]= 1197050035;
assign addr[31064]= 1259782632;
assign addr[31065]= 1320917099;
assign addr[31066]= 1380375881;
assign addr[31067]= 1438083551;
assign addr[31068]= 1493966902;
assign addr[31069]= 1547955041;
assign addr[31070]= 1599979481;
assign addr[31071]= 1649974225;
assign addr[31072]= 1697875851;
assign addr[31073]= 1743623590;
assign addr[31074]= 1787159411;
assign addr[31075]= 1828428082;
assign addr[31076]= 1867377253;
assign addr[31077]= 1903957513;
assign addr[31078]= 1938122457;
assign addr[31079]= 1969828744;
assign addr[31080]= 1999036154;
assign addr[31081]= 2025707632;
assign addr[31082]= 2049809346;
assign addr[31083]= 2071310720;
assign addr[31084]= 2090184478;
assign addr[31085]= 2106406677;
assign addr[31086]= 2119956737;
assign addr[31087]= 2130817471;
assign addr[31088]= 2138975100;
assign addr[31089]= 2144419275;
assign addr[31090]= 2147143090;
assign addr[31091]= 2147143090;
assign addr[31092]= 2144419275;
assign addr[31093]= 2138975100;
assign addr[31094]= 2130817471;
assign addr[31095]= 2119956737;
assign addr[31096]= 2106406677;
assign addr[31097]= 2090184478;
assign addr[31098]= 2071310720;
assign addr[31099]= 2049809346;
assign addr[31100]= 2025707632;
assign addr[31101]= 1999036154;
assign addr[31102]= 1969828744;
assign addr[31103]= 1938122457;
assign addr[31104]= 1903957513;
assign addr[31105]= 1867377253;
assign addr[31106]= 1828428082;
assign addr[31107]= 1787159411;
assign addr[31108]= 1743623590;
assign addr[31109]= 1697875851;
assign addr[31110]= 1649974225;
assign addr[31111]= 1599979481;
assign addr[31112]= 1547955041;
assign addr[31113]= 1493966902;
assign addr[31114]= 1438083551;
assign addr[31115]= 1380375881;
assign addr[31116]= 1320917099;
assign addr[31117]= 1259782632;
assign addr[31118]= 1197050035;
assign addr[31119]= 1132798888;
assign addr[31120]= 1067110699;
assign addr[31121]= 1000068799;
assign addr[31122]= 931758235;
assign addr[31123]= 862265664;
assign addr[31124]= 791679244;
assign addr[31125]= 720088517;
assign addr[31126]= 647584304;
assign addr[31127]= 574258580;
assign addr[31128]= 500204365;
assign addr[31129]= 425515602;
assign addr[31130]= 350287041;
assign addr[31131]= 274614114;
assign addr[31132]= 198592817;
assign addr[31133]= 122319591;
assign addr[31134]= 45891193;
assign addr[31135]= -30595422;
assign addr[31136]= -107043224;
assign addr[31137]= -183355234;
assign addr[31138]= -259434643;
assign addr[31139]= -335184940;
assign addr[31140]= -410510029;
assign addr[31141]= -485314355;
assign addr[31142]= -559503022;
assign addr[31143]= -632981917;
assign addr[31144]= -705657826;
assign addr[31145]= -777438554;
assign addr[31146]= -848233042;
assign addr[31147]= -917951481;
assign addr[31148]= -986505429;
assign addr[31149]= -1053807919;
assign addr[31150]= -1119773573;
assign addr[31151]= -1184318708;
assign addr[31152]= -1247361445;
assign addr[31153]= -1308821808;
assign addr[31154]= -1368621831;
assign addr[31155]= -1426685652;
assign addr[31156]= -1482939614;
assign addr[31157]= -1537312353;
assign addr[31158]= -1589734894;
assign addr[31159]= -1640140734;
assign addr[31160]= -1688465931;
assign addr[31161]= -1734649179;
assign addr[31162]= -1778631892;
assign addr[31163]= -1820358275;
assign addr[31164]= -1859775393;
assign addr[31165]= -1896833245;
assign addr[31166]= -1931484818;
assign addr[31167]= -1963686155;
assign addr[31168]= -1993396407;
assign addr[31169]= -2020577882;
assign addr[31170]= -2045196100;
assign addr[31171]= -2067219829;
assign addr[31172]= -2086621133;
assign addr[31173]= -2103375398;
assign addr[31174]= -2117461370;
assign addr[31175]= -2128861181;
assign addr[31176]= -2137560369;
assign addr[31177]= -2143547897;
assign addr[31178]= -2146816171;
assign addr[31179]= -2147361045;
assign addr[31180]= -2145181827;
assign addr[31181]= -2140281282;
assign addr[31182]= -2132665626;
assign addr[31183]= -2122344521;
assign addr[31184]= -2109331059;
assign addr[31185]= -2093641749;
assign addr[31186]= -2075296495;
assign addr[31187]= -2054318569;
assign addr[31188]= -2030734582;
assign addr[31189]= -2004574453;
assign addr[31190]= -1975871368;
assign addr[31191]= -1944661739;
assign addr[31192]= -1910985158;
assign addr[31193]= -1874884346;
assign addr[31194]= -1836405100;
assign addr[31195]= -1795596234;
assign addr[31196]= -1752509516;
assign addr[31197]= -1707199606;
assign addr[31198]= -1659723983;
assign addr[31199]= -1610142873;
assign addr[31200]= -1558519173;
assign addr[31201]= -1504918373;
assign addr[31202]= -1449408469;
assign addr[31203]= -1392059879;
assign addr[31204]= -1332945355;
assign addr[31205]= -1272139887;
assign addr[31206]= -1209720613;
assign addr[31207]= -1145766716;
assign addr[31208]= -1080359326;
assign addr[31209]= -1013581418;
assign addr[31210]= -945517704;
assign addr[31211]= -876254528;
assign addr[31212]= -805879757;
assign addr[31213]= -734482665;
assign addr[31214]= -662153826;
assign addr[31215]= -588984994;
assign addr[31216]= -515068990;
assign addr[31217]= -440499581;
assign addr[31218]= -365371365;
assign addr[31219]= -289779648;
assign addr[31220]= -213820322;
assign addr[31221]= -137589750;
assign addr[31222]= -61184634;
assign addr[31223]= 15298099;
assign addr[31224]= 91761426;
assign addr[31225]= 168108346;
assign addr[31226]= 244242007;
assign addr[31227]= 320065829;
assign addr[31228]= 395483624;
assign addr[31229]= 470399716;
assign addr[31230]= 544719071;
assign addr[31231]= 618347408;
assign addr[31232]= 691191324;
assign addr[31233]= 763158411;
assign addr[31234]= 834157373;
assign addr[31235]= 904098143;
assign addr[31236]= 972891995;
assign addr[31237]= 1040451659;
assign addr[31238]= 1106691431;
assign addr[31239]= 1171527280;
assign addr[31240]= 1234876957;
assign addr[31241]= 1296660098;
assign addr[31242]= 1356798326;
assign addr[31243]= 1415215352;
assign addr[31244]= 1471837070;
assign addr[31245]= 1526591649;
assign addr[31246]= 1579409630;
assign addr[31247]= 1630224009;
assign addr[31248]= 1678970324;
assign addr[31249]= 1725586737;
assign addr[31250]= 1770014111;
assign addr[31251]= 1812196087;
assign addr[31252]= 1852079154;
assign addr[31253]= 1889612716;
assign addr[31254]= 1924749160;
assign addr[31255]= 1957443913;
assign addr[31256]= 1987655498;
assign addr[31257]= 2015345591;
assign addr[31258]= 2040479063;
assign addr[31259]= 2063024031;
assign addr[31260]= 2082951896;
assign addr[31261]= 2100237377;
assign addr[31262]= 2114858546;
assign addr[31263]= 2126796855;
assign addr[31264]= 2136037160;
assign addr[31265]= 2142567738;
assign addr[31266]= 2146380306;
assign addr[31267]= 2147470025;
assign addr[31268]= 2145835515;
assign addr[31269]= 2141478848;
assign addr[31270]= 2134405552;
assign addr[31271]= 2124624598;
assign addr[31272]= 2112148396;
assign addr[31273]= 2096992772;
assign addr[31274]= 2079176953;
assign addr[31275]= 2058723538;
assign addr[31276]= 2035658475;
assign addr[31277]= 2010011024;
assign addr[31278]= 1981813720;
assign addr[31279]= 1951102334;
assign addr[31280]= 1917915825;
assign addr[31281]= 1882296293;
assign addr[31282]= 1844288924;
assign addr[31283]= 1803941934;
assign addr[31284]= 1761306505;
assign addr[31285]= 1716436725;
assign addr[31286]= 1669389513;
assign addr[31287]= 1620224553;
assign addr[31288]= 1569004214;
assign addr[31289]= 1515793473;
assign addr[31290]= 1460659832;
assign addr[31291]= 1403673233;
assign addr[31292]= 1344905966;
assign addr[31293]= 1284432584;
assign addr[31294]= 1222329801;
assign addr[31295]= 1158676398;
assign addr[31296]= 1093553126;
assign addr[31297]= 1027042599;
assign addr[31298]= 959229189;
assign addr[31299]= 890198924;
assign addr[31300]= 820039373;
assign addr[31301]= 748839539;
assign addr[31302]= 676689746;
assign addr[31303]= 603681519;
assign addr[31304]= 529907477;
assign addr[31305]= 455461206;
assign addr[31306]= 380437148;
assign addr[31307]= 304930476;
assign addr[31308]= 229036977;
assign addr[31309]= 152852926;
assign addr[31310]= 76474970;
assign addr[31311]= 0;
assign addr[31312]= -76474970;
assign addr[31313]= -152852926;
assign addr[31314]= -229036977;
assign addr[31315]= -304930476;
assign addr[31316]= -380437148;
assign addr[31317]= -455461206;
assign addr[31318]= -529907477;
assign addr[31319]= -603681519;
assign addr[31320]= -676689746;
assign addr[31321]= -748839539;
assign addr[31322]= -820039373;
assign addr[31323]= -890198924;
assign addr[31324]= -959229189;
assign addr[31325]= -1027042599;
assign addr[31326]= -1093553126;
assign addr[31327]= -1158676398;
assign addr[31328]= -1222329801;
assign addr[31329]= -1284432584;
assign addr[31330]= -1344905966;
assign addr[31331]= -1403673233;
assign addr[31332]= -1460659832;
assign addr[31333]= -1515793473;
assign addr[31334]= -1569004214;
assign addr[31335]= -1620224553;
assign addr[31336]= -1669389513;
assign addr[31337]= -1716436725;
assign addr[31338]= -1761306505;
assign addr[31339]= -1803941934;
assign addr[31340]= -1844288924;
assign addr[31341]= -1882296293;
assign addr[31342]= -1917915825;
assign addr[31343]= -1951102334;
assign addr[31344]= -1981813720;
assign addr[31345]= -2010011024;
assign addr[31346]= -2035658475;
assign addr[31347]= -2058723538;
assign addr[31348]= -2079176953;
assign addr[31349]= -2096992772;
assign addr[31350]= -2112148396;
assign addr[31351]= -2124624598;
assign addr[31352]= -2134405552;
assign addr[31353]= -2141478848;
assign addr[31354]= -2145835515;
assign addr[31355]= -2147470025;
assign addr[31356]= -2146380306;
assign addr[31357]= -2142567738;
assign addr[31358]= -2136037160;
assign addr[31359]= -2126796855;
assign addr[31360]= -2114858546;
assign addr[31361]= -2100237377;
assign addr[31362]= -2082951896;
assign addr[31363]= -2063024031;
assign addr[31364]= -2040479063;
assign addr[31365]= -2015345591;
assign addr[31366]= -1987655498;
assign addr[31367]= -1957443913;
assign addr[31368]= -1924749160;
assign addr[31369]= -1889612716;
assign addr[31370]= -1852079154;
assign addr[31371]= -1812196087;
assign addr[31372]= -1770014111;
assign addr[31373]= -1725586737;
assign addr[31374]= -1678970324;
assign addr[31375]= -1630224009;
assign addr[31376]= -1579409630;
assign addr[31377]= -1526591649;
assign addr[31378]= -1471837070;
assign addr[31379]= -1415215352;
assign addr[31380]= -1356798326;
assign addr[31381]= -1296660098;
assign addr[31382]= -1234876957;
assign addr[31383]= -1171527280;
assign addr[31384]= -1106691431;
assign addr[31385]= -1040451659;
assign addr[31386]= -972891995;
assign addr[31387]= -904098143;
assign addr[31388]= -834157373;
assign addr[31389]= -763158411;
assign addr[31390]= -691191324;
assign addr[31391]= -618347408;
assign addr[31392]= -544719071;
assign addr[31393]= -470399716;
assign addr[31394]= -395483624;
assign addr[31395]= -320065829;
assign addr[31396]= -244242007;
assign addr[31397]= -168108346;
assign addr[31398]= -91761426;
assign addr[31399]= -15298099;
assign addr[31400]= 61184634;
assign addr[31401]= 137589750;
assign addr[31402]= 213820322;
assign addr[31403]= 289779648;
assign addr[31404]= 365371365;
assign addr[31405]= 440499581;
assign addr[31406]= 515068990;
assign addr[31407]= 588984994;
assign addr[31408]= 662153826;
assign addr[31409]= 734482665;
assign addr[31410]= 805879757;
assign addr[31411]= 876254528;
assign addr[31412]= 945517704;
assign addr[31413]= 1013581418;
assign addr[31414]= 1080359326;
assign addr[31415]= 1145766716;
assign addr[31416]= 1209720613;
assign addr[31417]= 1272139887;
assign addr[31418]= 1332945355;
assign addr[31419]= 1392059879;
assign addr[31420]= 1449408469;
assign addr[31421]= 1504918373;
assign addr[31422]= 1558519173;
assign addr[31423]= 1610142873;
assign addr[31424]= 1659723983;
assign addr[31425]= 1707199606;
assign addr[31426]= 1752509516;
assign addr[31427]= 1795596234;
assign addr[31428]= 1836405100;
assign addr[31429]= 1874884346;
assign addr[31430]= 1910985158;
assign addr[31431]= 1944661739;
assign addr[31432]= 1975871368;
assign addr[31433]= 2004574453;
assign addr[31434]= 2030734582;
assign addr[31435]= 2054318569;
assign addr[31436]= 2075296495;
assign addr[31437]= 2093641749;
assign addr[31438]= 2109331059;
assign addr[31439]= 2122344521;
assign addr[31440]= 2132665626;
assign addr[31441]= 2140281282;
assign addr[31442]= 2145181827;
assign addr[31443]= 2147361045;
assign addr[31444]= 2146816171;
assign addr[31445]= 2143547897;
assign addr[31446]= 2137560369;
assign addr[31447]= 2128861181;
assign addr[31448]= 2117461370;
assign addr[31449]= 2103375398;
assign addr[31450]= 2086621133;
assign addr[31451]= 2067219829;
assign addr[31452]= 2045196100;
assign addr[31453]= 2020577882;
assign addr[31454]= 1993396407;
assign addr[31455]= 1963686155;
assign addr[31456]= 1931484818;
assign addr[31457]= 1896833245;
assign addr[31458]= 1859775393;
assign addr[31459]= 1820358275;
assign addr[31460]= 1778631892;
assign addr[31461]= 1734649179;
assign addr[31462]= 1688465931;
assign addr[31463]= 1640140734;
assign addr[31464]= 1589734894;
assign addr[31465]= 1537312353;
assign addr[31466]= 1482939614;
assign addr[31467]= 1426685652;
assign addr[31468]= 1368621831;
assign addr[31469]= 1308821808;
assign addr[31470]= 1247361445;
assign addr[31471]= 1184318708;
assign addr[31472]= 1119773573;
assign addr[31473]= 1053807919;
assign addr[31474]= 986505429;
assign addr[31475]= 917951481;
assign addr[31476]= 848233042;
assign addr[31477]= 777438554;
assign addr[31478]= 705657826;
assign addr[31479]= 632981917;
assign addr[31480]= 559503022;
assign addr[31481]= 485314355;
assign addr[31482]= 410510029;
assign addr[31483]= 335184940;
assign addr[31484]= 259434643;
assign addr[31485]= 183355234;
assign addr[31486]= 107043224;
assign addr[31487]= 30595422;
assign addr[31488]= -45891193;
assign addr[31489]= -122319591;
assign addr[31490]= -198592817;
assign addr[31491]= -274614114;
assign addr[31492]= -350287041;
assign addr[31493]= -425515602;
assign addr[31494]= -500204365;
assign addr[31495]= -574258580;
assign addr[31496]= -647584304;
assign addr[31497]= -720088517;
assign addr[31498]= -791679244;
assign addr[31499]= -862265664;
assign addr[31500]= -931758235;
assign addr[31501]= -1000068799;
assign addr[31502]= -1067110699;
assign addr[31503]= -1132798888;
assign addr[31504]= -1197050035;
assign addr[31505]= -1259782632;
assign addr[31506]= -1320917099;
assign addr[31507]= -1380375881;
assign addr[31508]= -1438083551;
assign addr[31509]= -1493966902;
assign addr[31510]= -1547955041;
assign addr[31511]= -1599979481;
assign addr[31512]= -1649974225;
assign addr[31513]= -1697875851;
assign addr[31514]= -1743623590;
assign addr[31515]= -1787159411;
assign addr[31516]= -1828428082;
assign addr[31517]= -1867377253;
assign addr[31518]= -1903957513;
assign addr[31519]= -1938122457;
assign addr[31520]= -1969828744;
assign addr[31521]= -1999036154;
assign addr[31522]= -2025707632;
assign addr[31523]= -2049809346;
assign addr[31524]= -2071310720;
assign addr[31525]= -2090184478;
assign addr[31526]= -2106406677;
assign addr[31527]= -2119956737;
assign addr[31528]= -2130817471;
assign addr[31529]= -2138975100;
assign addr[31530]= -2144419275;
assign addr[31531]= -2147143090;
assign addr[31532]= -2147143090;
assign addr[31533]= -2144419275;
assign addr[31534]= -2138975100;
assign addr[31535]= -2130817471;
assign addr[31536]= -2119956737;
assign addr[31537]= -2106406677;
assign addr[31538]= -2090184478;
assign addr[31539]= -2071310720;
assign addr[31540]= -2049809346;
assign addr[31541]= -2025707632;
assign addr[31542]= -1999036154;
assign addr[31543]= -1969828744;
assign addr[31544]= -1938122457;
assign addr[31545]= -1903957513;
assign addr[31546]= -1867377253;
assign addr[31547]= -1828428082;
assign addr[31548]= -1787159411;
assign addr[31549]= -1743623590;
assign addr[31550]= -1697875851;
assign addr[31551]= -1649974225;
assign addr[31552]= -1599979481;
assign addr[31553]= -1547955041;
assign addr[31554]= -1493966902;
assign addr[31555]= -1438083551;
assign addr[31556]= -1380375881;
assign addr[31557]= -1320917099;
assign addr[31558]= -1259782632;
assign addr[31559]= -1197050035;
assign addr[31560]= -1132798888;
assign addr[31561]= -1067110699;
assign addr[31562]= -1000068799;
assign addr[31563]= -931758235;
assign addr[31564]= -862265664;
assign addr[31565]= -791679244;
assign addr[31566]= -720088517;
assign addr[31567]= -647584304;
assign addr[31568]= -574258580;
assign addr[31569]= -500204365;
assign addr[31570]= -425515602;
assign addr[31571]= -350287041;
assign addr[31572]= -274614114;
assign addr[31573]= -198592817;
assign addr[31574]= -122319591;
assign addr[31575]= -45891193;
assign addr[31576]= 30595422;
assign addr[31577]= 107043224;
assign addr[31578]= 183355234;
assign addr[31579]= 259434643;
assign addr[31580]= 335184940;
assign addr[31581]= 410510029;
assign addr[31582]= 485314355;
assign addr[31583]= 559503022;
assign addr[31584]= 632981917;
assign addr[31585]= 705657826;
assign addr[31586]= 777438554;
assign addr[31587]= 848233042;
assign addr[31588]= 917951481;
assign addr[31589]= 986505429;
assign addr[31590]= 1053807919;
assign addr[31591]= 1119773573;
assign addr[31592]= 1184318708;
assign addr[31593]= 1247361445;
assign addr[31594]= 1308821808;
assign addr[31595]= 1368621831;
assign addr[31596]= 1426685652;
assign addr[31597]= 1482939614;
assign addr[31598]= 1537312353;
assign addr[31599]= 1589734894;
assign addr[31600]= 1640140734;
assign addr[31601]= 1688465931;
assign addr[31602]= 1734649179;
assign addr[31603]= 1778631892;
assign addr[31604]= 1820358275;
assign addr[31605]= 1859775393;
assign addr[31606]= 1896833245;
assign addr[31607]= 1931484818;
assign addr[31608]= 1963686155;
assign addr[31609]= 1993396407;
assign addr[31610]= 2020577882;
assign addr[31611]= 2045196100;
assign addr[31612]= 2067219829;
assign addr[31613]= 2086621133;
assign addr[31614]= 2103375398;
assign addr[31615]= 2117461370;
assign addr[31616]= 2128861181;
assign addr[31617]= 2137560369;
assign addr[31618]= 2143547897;
assign addr[31619]= 2146816171;
assign addr[31620]= 2147361045;
assign addr[31621]= 2145181827;
assign addr[31622]= 2140281282;
assign addr[31623]= 2132665626;
assign addr[31624]= 2122344521;
assign addr[31625]= 2109331059;
assign addr[31626]= 2093641749;
assign addr[31627]= 2075296495;
assign addr[31628]= 2054318569;
assign addr[31629]= 2030734582;
assign addr[31630]= 2004574453;
assign addr[31631]= 1975871368;
assign addr[31632]= 1944661739;
assign addr[31633]= 1910985158;
assign addr[31634]= 1874884346;
assign addr[31635]= 1836405100;
assign addr[31636]= 1795596234;
assign addr[31637]= 1752509516;
assign addr[31638]= 1707199606;
assign addr[31639]= 1659723983;
assign addr[31640]= 1610142873;
assign addr[31641]= 1558519173;
assign addr[31642]= 1504918373;
assign addr[31643]= 1449408469;
assign addr[31644]= 1392059879;
assign addr[31645]= 1332945355;
assign addr[31646]= 1272139887;
assign addr[31647]= 1209720613;
assign addr[31648]= 1145766716;
assign addr[31649]= 1080359326;
assign addr[31650]= 1013581418;
assign addr[31651]= 945517704;
assign addr[31652]= 876254528;
assign addr[31653]= 805879757;
assign addr[31654]= 734482665;
assign addr[31655]= 662153826;
assign addr[31656]= 588984994;
assign addr[31657]= 515068990;
assign addr[31658]= 440499581;
assign addr[31659]= 365371365;
assign addr[31660]= 289779648;
assign addr[31661]= 213820322;
assign addr[31662]= 137589750;
assign addr[31663]= 61184634;
assign addr[31664]= -15298099;
assign addr[31665]= -91761426;
assign addr[31666]= -168108346;
assign addr[31667]= -244242007;
assign addr[31668]= -320065829;
assign addr[31669]= -395483624;
assign addr[31670]= -470399716;
assign addr[31671]= -544719071;
assign addr[31672]= -618347408;
assign addr[31673]= -691191324;
assign addr[31674]= -763158411;
assign addr[31675]= -834157373;
assign addr[31676]= -904098143;
assign addr[31677]= -972891995;
assign addr[31678]= -1040451659;
assign addr[31679]= -1106691431;
assign addr[31680]= -1171527280;
assign addr[31681]= -1234876957;
assign addr[31682]= -1296660098;
assign addr[31683]= -1356798326;
assign addr[31684]= -1415215352;
assign addr[31685]= -1471837070;
assign addr[31686]= -1526591649;
assign addr[31687]= -1579409630;
assign addr[31688]= -1630224009;
assign addr[31689]= -1678970324;
assign addr[31690]= -1725586737;
assign addr[31691]= -1770014111;
assign addr[31692]= -1812196087;
assign addr[31693]= -1852079154;
assign addr[31694]= -1889612716;
assign addr[31695]= -1924749160;
assign addr[31696]= -1957443913;
assign addr[31697]= -1987655498;
assign addr[31698]= -2015345591;
assign addr[31699]= -2040479063;
assign addr[31700]= -2063024031;
assign addr[31701]= -2082951896;
assign addr[31702]= -2100237377;
assign addr[31703]= -2114858546;
assign addr[31704]= -2126796855;
assign addr[31705]= -2136037160;
assign addr[31706]= -2142567738;
assign addr[31707]= -2146380306;
assign addr[31708]= -2147470025;
assign addr[31709]= -2145835515;
assign addr[31710]= -2141478848;
assign addr[31711]= -2134405552;
assign addr[31712]= -2124624598;
assign addr[31713]= -2112148396;
assign addr[31714]= -2096992772;
assign addr[31715]= -2079176953;
assign addr[31716]= -2058723538;
assign addr[31717]= -2035658475;
assign addr[31718]= -2010011024;
assign addr[31719]= -1981813720;
assign addr[31720]= -1951102334;
assign addr[31721]= -1917915825;
assign addr[31722]= -1882296293;
assign addr[31723]= -1844288924;
assign addr[31724]= -1803941934;
assign addr[31725]= -1761306505;
assign addr[31726]= -1716436725;
assign addr[31727]= -1669389513;
assign addr[31728]= -1620224553;
assign addr[31729]= -1569004214;
assign addr[31730]= -1515793473;
assign addr[31731]= -1460659832;
assign addr[31732]= -1403673233;
assign addr[31733]= -1344905966;
assign addr[31734]= -1284432584;
assign addr[31735]= -1222329801;
assign addr[31736]= -1158676398;
assign addr[31737]= -1093553126;
assign addr[31738]= -1027042599;
assign addr[31739]= -959229189;
assign addr[31740]= -890198924;
assign addr[31741]= -820039373;
assign addr[31742]= -748839539;
assign addr[31743]= -676689746;
assign addr[31744]= -603681519;
assign addr[31745]= -529907477;
assign addr[31746]= -455461206;
assign addr[31747]= -380437148;
assign addr[31748]= -304930476;
assign addr[31749]= -229036977;
assign addr[31750]= -152852926;
assign addr[31751]= -76474970;
assign addr[31752]= 0;
assign addr[31753]= 76474970;
assign addr[31754]= 152852926;
assign addr[31755]= 229036977;
assign addr[31756]= 304930476;
assign addr[31757]= 380437148;
assign addr[31758]= 455461206;
assign addr[31759]= 529907477;
assign addr[31760]= 603681519;
assign addr[31761]= 676689746;
assign addr[31762]= 748839539;
assign addr[31763]= 820039373;
assign addr[31764]= 890198924;
assign addr[31765]= 959229189;
assign addr[31766]= 1027042599;
assign addr[31767]= 1093553126;
assign addr[31768]= 1158676398;
assign addr[31769]= 1222329801;
assign addr[31770]= 1284432584;
assign addr[31771]= 1344905966;
assign addr[31772]= 1403673233;
assign addr[31773]= 1460659832;
assign addr[31774]= 1515793473;
assign addr[31775]= 1569004214;
assign addr[31776]= 1620224553;
assign addr[31777]= 1669389513;
assign addr[31778]= 1716436725;
assign addr[31779]= 1761306505;
assign addr[31780]= 1803941934;
assign addr[31781]= 1844288924;
assign addr[31782]= 1882296293;
assign addr[31783]= 1917915825;
assign addr[31784]= 1951102334;
assign addr[31785]= 1981813720;
assign addr[31786]= 2010011024;
assign addr[31787]= 2035658475;
assign addr[31788]= 2058723538;
assign addr[31789]= 2079176953;
assign addr[31790]= 2096992772;
assign addr[31791]= 2112148396;
assign addr[31792]= 2124624598;
assign addr[31793]= 2134405552;
assign addr[31794]= 2141478848;
assign addr[31795]= 2145835515;
assign addr[31796]= 2147470025;
assign addr[31797]= 2146380306;
assign addr[31798]= 2142567738;
assign addr[31799]= 2136037160;
assign addr[31800]= 2126796855;
assign addr[31801]= 2114858546;
assign addr[31802]= 2100237377;
assign addr[31803]= 2082951896;
assign addr[31804]= 2063024031;
assign addr[31805]= 2040479063;
assign addr[31806]= 2015345591;
assign addr[31807]= 1987655498;
assign addr[31808]= 1957443913;
assign addr[31809]= 1924749160;
assign addr[31810]= 1889612716;
assign addr[31811]= 1852079154;
assign addr[31812]= 1812196087;
assign addr[31813]= 1770014111;
assign addr[31814]= 1725586737;
assign addr[31815]= 1678970324;
assign addr[31816]= 1630224009;
assign addr[31817]= 1579409630;
assign addr[31818]= 1526591649;
assign addr[31819]= 1471837070;
assign addr[31820]= 1415215352;
assign addr[31821]= 1356798326;
assign addr[31822]= 1296660098;
assign addr[31823]= 1234876957;
assign addr[31824]= 1171527280;
assign addr[31825]= 1106691431;
assign addr[31826]= 1040451659;
assign addr[31827]= 972891995;
assign addr[31828]= 904098143;
assign addr[31829]= 834157373;
assign addr[31830]= 763158411;
assign addr[31831]= 691191324;
assign addr[31832]= 618347408;
assign addr[31833]= 544719071;
assign addr[31834]= 470399716;
assign addr[31835]= 395483624;
assign addr[31836]= 320065829;
assign addr[31837]= 244242007;
assign addr[31838]= 168108346;
assign addr[31839]= 91761426;
assign addr[31840]= 15298099;
assign addr[31841]= -61184634;
assign addr[31842]= -137589750;
assign addr[31843]= -213820322;
assign addr[31844]= -289779648;
assign addr[31845]= -365371365;
assign addr[31846]= -440499581;
assign addr[31847]= -515068990;
assign addr[31848]= -588984994;
assign addr[31849]= -662153826;
assign addr[31850]= -734482665;
assign addr[31851]= -805879757;
assign addr[31852]= -876254528;
assign addr[31853]= -945517704;
assign addr[31854]= -1013581418;
assign addr[31855]= -1080359326;
assign addr[31856]= -1145766716;
assign addr[31857]= -1209720613;
assign addr[31858]= -1272139887;
assign addr[31859]= -1332945355;
assign addr[31860]= -1392059879;
assign addr[31861]= -1449408469;
assign addr[31862]= -1504918373;
assign addr[31863]= -1558519173;
assign addr[31864]= -1610142873;
assign addr[31865]= -1659723983;
assign addr[31866]= -1707199606;
assign addr[31867]= -1752509516;
assign addr[31868]= -1795596234;
assign addr[31869]= -1836405100;
assign addr[31870]= -1874884346;
assign addr[31871]= -1910985158;
assign addr[31872]= -1944661739;
assign addr[31873]= -1975871368;
assign addr[31874]= -2004574453;
assign addr[31875]= -2030734582;
assign addr[31876]= -2054318569;
assign addr[31877]= -2075296495;
assign addr[31878]= -2093641749;
assign addr[31879]= -2109331059;
assign addr[31880]= -2122344521;
assign addr[31881]= -2132665626;
assign addr[31882]= -2140281282;
assign addr[31883]= -2145181827;
assign addr[31884]= -2147361045;
assign addr[31885]= -2146816171;
assign addr[31886]= -2143547897;
assign addr[31887]= -2137560369;
assign addr[31888]= -2128861181;
assign addr[31889]= -2117461370;
assign addr[31890]= -2103375398;
assign addr[31891]= -2086621133;
assign addr[31892]= -2067219829;
assign addr[31893]= -2045196100;
assign addr[31894]= -2020577882;
assign addr[31895]= -1993396407;
assign addr[31896]= -1963686155;
assign addr[31897]= -1931484818;
assign addr[31898]= -1896833245;
assign addr[31899]= -1859775393;
assign addr[31900]= -1820358275;
assign addr[31901]= -1778631892;
assign addr[31902]= -1734649179;
assign addr[31903]= -1688465931;
assign addr[31904]= -1640140734;
assign addr[31905]= -1589734894;
assign addr[31906]= -1537312353;
assign addr[31907]= -1482939614;
assign addr[31908]= -1426685652;
assign addr[31909]= -1368621831;
assign addr[31910]= -1308821808;
assign addr[31911]= -1247361445;
assign addr[31912]= -1184318708;
assign addr[31913]= -1119773573;
assign addr[31914]= -1053807919;
assign addr[31915]= -986505429;
assign addr[31916]= -917951481;
assign addr[31917]= -848233042;
assign addr[31918]= -777438554;
assign addr[31919]= -705657826;
assign addr[31920]= -632981917;
assign addr[31921]= -559503022;
assign addr[31922]= -485314355;
assign addr[31923]= -410510029;
assign addr[31924]= -335184940;
assign addr[31925]= -259434643;
assign addr[31926]= -183355234;
assign addr[31927]= -107043224;
assign addr[31928]= -30595422;
assign addr[31929]= 45891193;
assign addr[31930]= 122319591;
assign addr[31931]= 198592817;
assign addr[31932]= 274614114;
assign addr[31933]= 350287041;
assign addr[31934]= 425515602;
assign addr[31935]= 500204365;
assign addr[31936]= 574258580;
assign addr[31937]= 647584304;
assign addr[31938]= 720088517;
assign addr[31939]= 791679244;
assign addr[31940]= 862265664;
assign addr[31941]= 931758235;
assign addr[31942]= 1000068799;
assign addr[31943]= 1067110699;
assign addr[31944]= 1132798888;
assign addr[31945]= 1197050035;
assign addr[31946]= 1259782632;
assign addr[31947]= 1320917099;
assign addr[31948]= 1380375881;
assign addr[31949]= 1438083551;
assign addr[31950]= 1493966902;
assign addr[31951]= 1547955041;
assign addr[31952]= 1599979481;
assign addr[31953]= 1649974225;
assign addr[31954]= 1697875851;
assign addr[31955]= 1743623590;
assign addr[31956]= 1787159411;
assign addr[31957]= 1828428082;
assign addr[31958]= 1867377253;
assign addr[31959]= 1903957513;
assign addr[31960]= 1938122457;
assign addr[31961]= 1969828744;
assign addr[31962]= 1999036154;
assign addr[31963]= 2025707632;
assign addr[31964]= 2049809346;
assign addr[31965]= 2071310720;
assign addr[31966]= 2090184478;
assign addr[31967]= 2106406677;
assign addr[31968]= 2119956737;
assign addr[31969]= 2130817471;
assign addr[31970]= 2138975100;
assign addr[31971]= 2144419275;
assign addr[31972]= 2147143090;
assign addr[31973]= 2147143090;
assign addr[31974]= 2144419275;
assign addr[31975]= 2138975100;
assign addr[31976]= 2130817471;
assign addr[31977]= 2119956737;
assign addr[31978]= 2106406677;
assign addr[31979]= 2090184478;
assign addr[31980]= 2071310720;
assign addr[31981]= 2049809346;
assign addr[31982]= 2025707632;
assign addr[31983]= 1999036154;
assign addr[31984]= 1969828744;
assign addr[31985]= 1938122457;
assign addr[31986]= 1903957513;
assign addr[31987]= 1867377253;
assign addr[31988]= 1828428082;
assign addr[31989]= 1787159411;
assign addr[31990]= 1743623590;
assign addr[31991]= 1697875851;
assign addr[31992]= 1649974225;
assign addr[31993]= 1599979481;
assign addr[31994]= 1547955041;
assign addr[31995]= 1493966902;
assign addr[31996]= 1438083551;
assign addr[31997]= 1380375881;
assign addr[31998]= 1320917099;
assign addr[31999]= 1259782632;
assign addr[32000]= 1197050035;
assign addr[32001]= 1132798888;
assign addr[32002]= 1067110699;
assign addr[32003]= 1000068799;
assign addr[32004]= 931758235;
assign addr[32005]= 862265664;
assign addr[32006]= 791679244;
assign addr[32007]= 720088517;
assign addr[32008]= 647584304;
assign addr[32009]= 574258580;
assign addr[32010]= 500204365;
assign addr[32011]= 425515602;
assign addr[32012]= 350287041;
assign addr[32013]= 274614114;
assign addr[32014]= 198592817;
assign addr[32015]= 122319591;
assign addr[32016]= 45891193;
assign addr[32017]= -30595422;
assign addr[32018]= -107043224;
assign addr[32019]= -183355234;
assign addr[32020]= -259434643;
assign addr[32021]= -335184940;
assign addr[32022]= -410510029;
assign addr[32023]= -485314355;
assign addr[32024]= -559503022;
assign addr[32025]= -632981917;
assign addr[32026]= -705657826;
assign addr[32027]= -777438554;
assign addr[32028]= -848233042;
assign addr[32029]= -917951481;
assign addr[32030]= -986505429;
assign addr[32031]= -1053807919;
assign addr[32032]= -1119773573;
assign addr[32033]= -1184318708;
assign addr[32034]= -1247361445;
assign addr[32035]= -1308821808;
assign addr[32036]= -1368621831;
assign addr[32037]= -1426685652;
assign addr[32038]= -1482939614;
assign addr[32039]= -1537312353;
assign addr[32040]= -1589734894;
assign addr[32041]= -1640140734;
assign addr[32042]= -1688465931;
assign addr[32043]= -1734649179;
assign addr[32044]= -1778631892;
assign addr[32045]= -1820358275;
assign addr[32046]= -1859775393;
assign addr[32047]= -1896833245;
assign addr[32048]= -1931484818;
assign addr[32049]= -1963686155;
assign addr[32050]= -1993396407;
assign addr[32051]= -2020577882;
assign addr[32052]= -2045196100;
assign addr[32053]= -2067219829;
assign addr[32054]= -2086621133;
assign addr[32055]= -2103375398;
assign addr[32056]= -2117461370;
assign addr[32057]= -2128861181;
assign addr[32058]= -2137560369;
assign addr[32059]= -2143547897;
assign addr[32060]= -2146816171;
assign addr[32061]= -2147361045;
assign addr[32062]= -2145181827;
assign addr[32063]= -2140281282;
assign addr[32064]= -2132665626;
assign addr[32065]= -2122344521;
assign addr[32066]= -2109331059;
assign addr[32067]= -2093641749;
assign addr[32068]= -2075296495;
assign addr[32069]= -2054318569;
assign addr[32070]= -2030734582;
assign addr[32071]= -2004574453;
assign addr[32072]= -1975871368;
assign addr[32073]= -1944661739;
assign addr[32074]= -1910985158;
assign addr[32075]= -1874884346;
assign addr[32076]= -1836405100;
assign addr[32077]= -1795596234;
assign addr[32078]= -1752509516;
assign addr[32079]= -1707199606;
assign addr[32080]= -1659723983;
assign addr[32081]= -1610142873;
assign addr[32082]= -1558519173;
assign addr[32083]= -1504918373;
assign addr[32084]= -1449408469;
assign addr[32085]= -1392059879;
assign addr[32086]= -1332945355;
assign addr[32087]= -1272139887;
assign addr[32088]= -1209720613;
assign addr[32089]= -1145766716;
assign addr[32090]= -1080359326;
assign addr[32091]= -1013581418;
assign addr[32092]= -945517704;
assign addr[32093]= -876254528;
assign addr[32094]= -805879757;
assign addr[32095]= -734482665;
assign addr[32096]= -662153826;
assign addr[32097]= -588984994;
assign addr[32098]= -515068990;
assign addr[32099]= -440499581;
assign addr[32100]= -365371365;
assign addr[32101]= -289779648;
assign addr[32102]= -213820322;
assign addr[32103]= -137589750;
assign addr[32104]= -61184634;
assign addr[32105]= 15298099;
assign addr[32106]= 91761426;
assign addr[32107]= 168108346;
assign addr[32108]= 244242007;
assign addr[32109]= 320065829;
assign addr[32110]= 395483624;
assign addr[32111]= 470399716;
assign addr[32112]= 544719071;
assign addr[32113]= 618347408;
assign addr[32114]= 691191324;
assign addr[32115]= 763158411;
assign addr[32116]= 834157373;
assign addr[32117]= 904098143;
assign addr[32118]= 972891995;
assign addr[32119]= 1040451659;
assign addr[32120]= 1106691431;
assign addr[32121]= 1171527280;
assign addr[32122]= 1234876957;
assign addr[32123]= 1296660098;
assign addr[32124]= 1356798326;
assign addr[32125]= 1415215352;
assign addr[32126]= 1471837070;
assign addr[32127]= 1526591649;
assign addr[32128]= 1579409630;
assign addr[32129]= 1630224009;
assign addr[32130]= 1678970324;
assign addr[32131]= 1725586737;
assign addr[32132]= 1770014111;
assign addr[32133]= 1812196087;
assign addr[32134]= 1852079154;
assign addr[32135]= 1889612716;
assign addr[32136]= 1924749160;
assign addr[32137]= 1957443913;
assign addr[32138]= 1987655498;
assign addr[32139]= 2015345591;
assign addr[32140]= 2040479063;
assign addr[32141]= 2063024031;
assign addr[32142]= 2082951896;
assign addr[32143]= 2100237377;
assign addr[32144]= 2114858546;
assign addr[32145]= 2126796855;
assign addr[32146]= 2136037160;
assign addr[32147]= 2142567738;
assign addr[32148]= 2146380306;
assign addr[32149]= 2147470025;
assign addr[32150]= 2145835515;
assign addr[32151]= 2141478848;
assign addr[32152]= 2134405552;
assign addr[32153]= 2124624598;
assign addr[32154]= 2112148396;
assign addr[32155]= 2096992772;
assign addr[32156]= 2079176953;
assign addr[32157]= 2058723538;
assign addr[32158]= 2035658475;
assign addr[32159]= 2010011024;
assign addr[32160]= 1981813720;
assign addr[32161]= 1951102334;
assign addr[32162]= 1917915825;
assign addr[32163]= 1882296293;
assign addr[32164]= 1844288924;
assign addr[32165]= 1803941934;
assign addr[32166]= 1761306505;
assign addr[32167]= 1716436725;
assign addr[32168]= 1669389513;
assign addr[32169]= 1620224553;
assign addr[32170]= 1569004214;
assign addr[32171]= 1515793473;
assign addr[32172]= 1460659832;
assign addr[32173]= 1403673233;
assign addr[32174]= 1344905966;
assign addr[32175]= 1284432584;
assign addr[32176]= 1222329801;
assign addr[32177]= 1158676398;
assign addr[32178]= 1093553126;
assign addr[32179]= 1027042599;
assign addr[32180]= 959229189;
assign addr[32181]= 890198924;
assign addr[32182]= 820039373;
assign addr[32183]= 748839539;
assign addr[32184]= 676689746;
assign addr[32185]= 603681519;
assign addr[32186]= 529907477;
assign addr[32187]= 455461206;
assign addr[32188]= 380437148;
assign addr[32189]= 304930476;
assign addr[32190]= 229036977;
assign addr[32191]= 152852926;
assign addr[32192]= 76474970;
assign addr[32193]= 0;
assign addr[32194]= -76474970;
assign addr[32195]= -152852926;
assign addr[32196]= -229036977;
assign addr[32197]= -304930476;
assign addr[32198]= -380437148;
assign addr[32199]= -455461206;
assign addr[32200]= -529907477;
assign addr[32201]= -603681519;
assign addr[32202]= -676689746;
assign addr[32203]= -748839539;
assign addr[32204]= -820039373;
assign addr[32205]= -890198924;
assign addr[32206]= -959229189;
assign addr[32207]= -1027042599;
assign addr[32208]= -1093553126;
assign addr[32209]= -1158676398;
assign addr[32210]= -1222329801;
assign addr[32211]= -1284432584;
assign addr[32212]= -1344905966;
assign addr[32213]= -1403673233;
assign addr[32214]= -1460659832;
assign addr[32215]= -1515793473;
assign addr[32216]= -1569004214;
assign addr[32217]= -1620224553;
assign addr[32218]= -1669389513;
assign addr[32219]= -1716436725;
assign addr[32220]= -1761306505;
assign addr[32221]= -1803941934;
assign addr[32222]= -1844288924;
assign addr[32223]= -1882296293;
assign addr[32224]= -1917915825;
assign addr[32225]= -1951102334;
assign addr[32226]= -1981813720;
assign addr[32227]= -2010011024;
assign addr[32228]= -2035658475;
assign addr[32229]= -2058723538;
assign addr[32230]= -2079176953;
assign addr[32231]= -2096992772;
assign addr[32232]= -2112148396;
assign addr[32233]= -2124624598;
assign addr[32234]= -2134405552;
assign addr[32235]= -2141478848;
assign addr[32236]= -2145835515;
assign addr[32237]= -2147470025;
assign addr[32238]= -2146380306;
assign addr[32239]= -2142567738;
assign addr[32240]= -2136037160;
assign addr[32241]= -2126796855;
assign addr[32242]= -2114858546;
assign addr[32243]= -2100237377;
assign addr[32244]= -2082951896;
assign addr[32245]= -2063024031;
assign addr[32246]= -2040479063;
assign addr[32247]= -2015345591;
assign addr[32248]= -1987655498;
assign addr[32249]= -1957443913;
assign addr[32250]= -1924749160;
assign addr[32251]= -1889612716;
assign addr[32252]= -1852079154;
assign addr[32253]= -1812196087;
assign addr[32254]= -1770014111;
assign addr[32255]= -1725586737;
assign addr[32256]= -1678970324;
assign addr[32257]= -1630224009;
assign addr[32258]= -1579409630;
assign addr[32259]= -1526591649;
assign addr[32260]= -1471837070;
assign addr[32261]= -1415215352;
assign addr[32262]= -1356798326;
assign addr[32263]= -1296660098;
assign addr[32264]= -1234876957;
assign addr[32265]= -1171527280;
assign addr[32266]= -1106691431;
assign addr[32267]= -1040451659;
assign addr[32268]= -972891995;
assign addr[32269]= -904098143;
assign addr[32270]= -834157373;
assign addr[32271]= -763158411;
assign addr[32272]= -691191324;
assign addr[32273]= -618347408;
assign addr[32274]= -544719071;
assign addr[32275]= -470399716;
assign addr[32276]= -395483624;
assign addr[32277]= -320065829;
assign addr[32278]= -244242007;
assign addr[32279]= -168108346;
assign addr[32280]= -91761426;
assign addr[32281]= -15298099;
assign addr[32282]= 61184634;
assign addr[32283]= 137589750;
assign addr[32284]= 213820322;
assign addr[32285]= 289779648;
assign addr[32286]= 365371365;
assign addr[32287]= 440499581;
assign addr[32288]= 515068990;
assign addr[32289]= 588984994;
assign addr[32290]= 662153826;
assign addr[32291]= 734482665;
assign addr[32292]= 805879757;
assign addr[32293]= 876254528;
assign addr[32294]= 945517704;
assign addr[32295]= 1013581418;
assign addr[32296]= 1080359326;
assign addr[32297]= 1145766716;
assign addr[32298]= 1209720613;
assign addr[32299]= 1272139887;
assign addr[32300]= 1332945355;
assign addr[32301]= 1392059879;
assign addr[32302]= 1449408469;
assign addr[32303]= 1504918373;
assign addr[32304]= 1558519173;
assign addr[32305]= 1610142873;
assign addr[32306]= 1659723983;
assign addr[32307]= 1707199606;
assign addr[32308]= 1752509516;
assign addr[32309]= 1795596234;
assign addr[32310]= 1836405100;
assign addr[32311]= 1874884346;
assign addr[32312]= 1910985158;
assign addr[32313]= 1944661739;
assign addr[32314]= 1975871368;
assign addr[32315]= 2004574453;
assign addr[32316]= 2030734582;
assign addr[32317]= 2054318569;
assign addr[32318]= 2075296495;
assign addr[32319]= 2093641749;
assign addr[32320]= 2109331059;
assign addr[32321]= 2122344521;
assign addr[32322]= 2132665626;
assign addr[32323]= 2140281282;
assign addr[32324]= 2145181827;
assign addr[32325]= 2147361045;
assign addr[32326]= 2146816171;
assign addr[32327]= 2143547897;
assign addr[32328]= 2137560369;
assign addr[32329]= 2128861181;
assign addr[32330]= 2117461370;
assign addr[32331]= 2103375398;
assign addr[32332]= 2086621133;
assign addr[32333]= 2067219829;
assign addr[32334]= 2045196100;
assign addr[32335]= 2020577882;
assign addr[32336]= 1993396407;
assign addr[32337]= 1963686155;
assign addr[32338]= 1931484818;
assign addr[32339]= 1896833245;
assign addr[32340]= 1859775393;
assign addr[32341]= 1820358275;
assign addr[32342]= 1778631892;
assign addr[32343]= 1734649179;
assign addr[32344]= 1688465931;
assign addr[32345]= 1640140734;
assign addr[32346]= 1589734894;
assign addr[32347]= 1537312353;
assign addr[32348]= 1482939614;
assign addr[32349]= 1426685652;
assign addr[32350]= 1368621831;
assign addr[32351]= 1308821808;
assign addr[32352]= 1247361445;
assign addr[32353]= 1184318708;
assign addr[32354]= 1119773573;
assign addr[32355]= 1053807919;
assign addr[32356]= 986505429;
assign addr[32357]= 917951481;
assign addr[32358]= 848233042;
assign addr[32359]= 777438554;
assign addr[32360]= 705657826;
assign addr[32361]= 632981917;
assign addr[32362]= 559503022;
assign addr[32363]= 485314355;
assign addr[32364]= 410510029;
assign addr[32365]= 335184940;
assign addr[32366]= 259434643;
assign addr[32367]= 183355234;
assign addr[32368]= 107043224;
assign addr[32369]= 30595422;
assign addr[32370]= -45891193;
assign addr[32371]= -122319591;
assign addr[32372]= -198592817;
assign addr[32373]= -274614114;
assign addr[32374]= -350287041;
assign addr[32375]= -425515602;
assign addr[32376]= -500204365;
assign addr[32377]= -574258580;
assign addr[32378]= -647584304;
assign addr[32379]= -720088517;
assign addr[32380]= -791679244;
assign addr[32381]= -862265664;
assign addr[32382]= -931758235;
assign addr[32383]= -1000068799;
assign addr[32384]= -1067110699;
assign addr[32385]= -1132798888;
assign addr[32386]= -1197050035;
assign addr[32387]= -1259782632;
assign addr[32388]= -1320917099;
assign addr[32389]= -1380375881;
assign addr[32390]= -1438083551;
assign addr[32391]= -1493966902;
assign addr[32392]= -1547955041;
assign addr[32393]= -1599979481;
assign addr[32394]= -1649974225;
assign addr[32395]= -1697875851;
assign addr[32396]= -1743623590;
assign addr[32397]= -1787159411;
assign addr[32398]= -1828428082;
assign addr[32399]= -1867377253;
assign addr[32400]= -1903957513;
assign addr[32401]= -1938122457;
assign addr[32402]= -1969828744;
assign addr[32403]= -1999036154;
assign addr[32404]= -2025707632;
assign addr[32405]= -2049809346;
assign addr[32406]= -2071310720;
assign addr[32407]= -2090184478;
assign addr[32408]= -2106406677;
assign addr[32409]= -2119956737;
assign addr[32410]= -2130817471;
assign addr[32411]= -2138975100;
assign addr[32412]= -2144419275;
assign addr[32413]= -2147143090;
assign addr[32414]= -2147143090;
assign addr[32415]= -2144419275;
assign addr[32416]= -2138975100;
assign addr[32417]= -2130817471;
assign addr[32418]= -2119956737;
assign addr[32419]= -2106406677;
assign addr[32420]= -2090184478;
assign addr[32421]= -2071310720;
assign addr[32422]= -2049809346;
assign addr[32423]= -2025707632;
assign addr[32424]= -1999036154;
assign addr[32425]= -1969828744;
assign addr[32426]= -1938122457;
assign addr[32427]= -1903957513;
assign addr[32428]= -1867377253;
assign addr[32429]= -1828428082;
assign addr[32430]= -1787159411;
assign addr[32431]= -1743623590;
assign addr[32432]= -1697875851;
assign addr[32433]= -1649974225;
assign addr[32434]= -1599979481;
assign addr[32435]= -1547955041;
assign addr[32436]= -1493966902;
assign addr[32437]= -1438083551;
assign addr[32438]= -1380375881;
assign addr[32439]= -1320917099;
assign addr[32440]= -1259782632;
assign addr[32441]= -1197050035;
assign addr[32442]= -1132798888;
assign addr[32443]= -1067110699;
assign addr[32444]= -1000068799;
assign addr[32445]= -931758235;
assign addr[32446]= -862265664;
assign addr[32447]= -791679244;
assign addr[32448]= -720088517;
assign addr[32449]= -647584304;
assign addr[32450]= -574258580;
assign addr[32451]= -500204365;
assign addr[32452]= -425515602;
assign addr[32453]= -350287041;
assign addr[32454]= -274614114;
assign addr[32455]= -198592817;
assign addr[32456]= -122319591;
assign addr[32457]= -45891193;
assign addr[32458]= 30595422;
assign addr[32459]= 107043224;
assign addr[32460]= 183355234;
assign addr[32461]= 259434643;
assign addr[32462]= 335184940;
assign addr[32463]= 410510029;
assign addr[32464]= 485314355;
assign addr[32465]= 559503022;
assign addr[32466]= 632981917;
assign addr[32467]= 705657826;
assign addr[32468]= 777438554;
assign addr[32469]= 848233042;
assign addr[32470]= 917951481;
assign addr[32471]= 986505429;
assign addr[32472]= 1053807919;
assign addr[32473]= 1119773573;
assign addr[32474]= 1184318708;
assign addr[32475]= 1247361445;
assign addr[32476]= 1308821808;
assign addr[32477]= 1368621831;
assign addr[32478]= 1426685652;
assign addr[32479]= 1482939614;
assign addr[32480]= 1537312353;
assign addr[32481]= 1589734894;
assign addr[32482]= 1640140734;
assign addr[32483]= 1688465931;
assign addr[32484]= 1734649179;
assign addr[32485]= 1778631892;
assign addr[32486]= 1820358275;
assign addr[32487]= 1859775393;
assign addr[32488]= 1896833245;
assign addr[32489]= 1931484818;
assign addr[32490]= 1963686155;
assign addr[32491]= 1993396407;
assign addr[32492]= 2020577882;
assign addr[32493]= 2045196100;
assign addr[32494]= 2067219829;
assign addr[32495]= 2086621133;
assign addr[32496]= 2103375398;
assign addr[32497]= 2117461370;
assign addr[32498]= 2128861181;
assign addr[32499]= 2137560369;
assign addr[32500]= 2143547897;
assign addr[32501]= 2146816171;
assign addr[32502]= 2147361045;
assign addr[32503]= 2145181827;
assign addr[32504]= 2140281282;
assign addr[32505]= 2132665626;
assign addr[32506]= 2122344521;
assign addr[32507]= 2109331059;
assign addr[32508]= 2093641749;
assign addr[32509]= 2075296495;
assign addr[32510]= 2054318569;
assign addr[32511]= 2030734582;
assign addr[32512]= 2004574453;
assign addr[32513]= 1975871368;
assign addr[32514]= 1944661739;
assign addr[32515]= 1910985158;
assign addr[32516]= 1874884346;
assign addr[32517]= 1836405100;
assign addr[32518]= 1795596234;
assign addr[32519]= 1752509516;
assign addr[32520]= 1707199606;
assign addr[32521]= 1659723983;
assign addr[32522]= 1610142873;
assign addr[32523]= 1558519173;
assign addr[32524]= 1504918373;
assign addr[32525]= 1449408469;
assign addr[32526]= 1392059879;
assign addr[32527]= 1332945355;
assign addr[32528]= 1272139887;
assign addr[32529]= 1209720613;
assign addr[32530]= 1145766716;
assign addr[32531]= 1080359326;
assign addr[32532]= 1013581418;
assign addr[32533]= 945517704;
assign addr[32534]= 876254528;
assign addr[32535]= 805879757;
assign addr[32536]= 734482665;
assign addr[32537]= 662153826;
assign addr[32538]= 588984994;
assign addr[32539]= 515068990;
assign addr[32540]= 440499581;
assign addr[32541]= 365371365;
assign addr[32542]= 289779648;
assign addr[32543]= 213820322;
assign addr[32544]= 137589750;
assign addr[32545]= 61184634;
assign addr[32546]= -15298099;
assign addr[32547]= -91761426;
assign addr[32548]= -168108346;
assign addr[32549]= -244242007;
assign addr[32550]= -320065829;
assign addr[32551]= -395483624;
assign addr[32552]= -470399716;
assign addr[32553]= -544719071;
assign addr[32554]= -618347408;
assign addr[32555]= -691191324;
assign addr[32556]= -763158411;
assign addr[32557]= -834157373;
assign addr[32558]= -904098143;
assign addr[32559]= -972891995;
assign addr[32560]= -1040451659;
assign addr[32561]= -1106691431;
assign addr[32562]= -1171527280;
assign addr[32563]= -1234876957;
assign addr[32564]= -1296660098;
assign addr[32565]= -1356798326;
assign addr[32566]= -1415215352;
assign addr[32567]= -1471837070;
assign addr[32568]= -1526591649;
assign addr[32569]= -1579409630;
assign addr[32570]= -1630224009;
assign addr[32571]= -1678970324;
assign addr[32572]= -1725586737;
assign addr[32573]= -1770014111;
assign addr[32574]= -1812196087;
assign addr[32575]= -1852079154;
assign addr[32576]= -1889612716;
assign addr[32577]= -1924749160;
assign addr[32578]= -1957443913;
assign addr[32579]= -1987655498;
assign addr[32580]= -2015345591;
assign addr[32581]= -2040479063;
assign addr[32582]= -2063024031;
assign addr[32583]= -2082951896;
assign addr[32584]= -2100237377;
assign addr[32585]= -2114858546;
assign addr[32586]= -2126796855;
assign addr[32587]= -2136037160;
assign addr[32588]= -2142567738;
assign addr[32589]= -2146380306;
assign addr[32590]= -2147470025;
assign addr[32591]= -2145835515;
assign addr[32592]= -2141478848;
assign addr[32593]= -2134405552;
assign addr[32594]= -2124624598;
assign addr[32595]= -2112148396;
assign addr[32596]= -2096992772;
assign addr[32597]= -2079176953;
assign addr[32598]= -2058723538;
assign addr[32599]= -2035658475;
assign addr[32600]= -2010011024;
assign addr[32601]= -1981813720;
assign addr[32602]= -1951102334;
assign addr[32603]= -1917915825;
assign addr[32604]= -1882296293;
assign addr[32605]= -1844288924;
assign addr[32606]= -1803941934;
assign addr[32607]= -1761306505;
assign addr[32608]= -1716436725;
assign addr[32609]= -1669389513;
assign addr[32610]= -1620224553;
assign addr[32611]= -1569004214;
assign addr[32612]= -1515793473;
assign addr[32613]= -1460659832;
assign addr[32614]= -1403673233;
assign addr[32615]= -1344905966;
assign addr[32616]= -1284432584;
assign addr[32617]= -1222329801;
assign addr[32618]= -1158676398;
assign addr[32619]= -1093553126;
assign addr[32620]= -1027042599;
assign addr[32621]= -959229189;
assign addr[32622]= -890198924;
assign addr[32623]= -820039373;
assign addr[32624]= -748839539;
assign addr[32625]= -676689746;
assign addr[32626]= -603681519;
assign addr[32627]= -529907477;
assign addr[32628]= -455461206;
assign addr[32629]= -380437148;
assign addr[32630]= -304930476;
assign addr[32631]= -229036977;
assign addr[32632]= -152852926;
assign addr[32633]= -76474970;
assign addr[32634]= 0;
assign addr[32635]= 76474970;
assign addr[32636]= 152852926;
assign addr[32637]= 229036977;
assign addr[32638]= 304930476;
assign addr[32639]= 380437148;
assign addr[32640]= 455461206;
assign addr[32641]= 529907477;
assign addr[32642]= 603681519;
assign addr[32643]= 676689746;
assign addr[32644]= 748839539;
assign addr[32645]= 820039373;
assign addr[32646]= 890198924;
assign addr[32647]= 959229189;
assign addr[32648]= 1027042599;
assign addr[32649]= 1093553126;
assign addr[32650]= 1158676398;
assign addr[32651]= 1222329801;
assign addr[32652]= 1284432584;
assign addr[32653]= 1344905966;
assign addr[32654]= 1403673233;
assign addr[32655]= 1460659832;
assign addr[32656]= 1515793473;
assign addr[32657]= 1569004214;
assign addr[32658]= 1620224553;
assign addr[32659]= 1669389513;
assign addr[32660]= 1716436725;
assign addr[32661]= 1761306505;
assign addr[32662]= 1803941934;
assign addr[32663]= 1844288924;
assign addr[32664]= 1882296293;
assign addr[32665]= 1917915825;
assign addr[32666]= 1951102334;
assign addr[32667]= 1981813720;
assign addr[32668]= 2010011024;
assign addr[32669]= 2035658475;
assign addr[32670]= 2058723538;
assign addr[32671]= 2079176953;
assign addr[32672]= 2096992772;
assign addr[32673]= 2112148396;
assign addr[32674]= 2124624598;
assign addr[32675]= 2134405552;
assign addr[32676]= 2141478848;
assign addr[32677]= 2145835515;
assign addr[32678]= 2147470025;
assign addr[32679]= 2146380306;
assign addr[32680]= 2142567738;
assign addr[32681]= 2136037160;
assign addr[32682]= 2126796855;
assign addr[32683]= 2114858546;
assign addr[32684]= 2100237377;
assign addr[32685]= 2082951896;
assign addr[32686]= 2063024031;
assign addr[32687]= 2040479063;
assign addr[32688]= 2015345591;
assign addr[32689]= 1987655498;
assign addr[32690]= 1957443913;
assign addr[32691]= 1924749160;
assign addr[32692]= 1889612716;
assign addr[32693]= 1852079154;
assign addr[32694]= 1812196087;
assign addr[32695]= 1770014111;
assign addr[32696]= 1725586737;
assign addr[32697]= 1678970324;
assign addr[32698]= 1630224009;
assign addr[32699]= 1579409630;
assign addr[32700]= 1526591649;
assign addr[32701]= 1471837070;
assign addr[32702]= 1415215352;
assign addr[32703]= 1356798326;
assign addr[32704]= 1296660098;
assign addr[32705]= 1234876957;
assign addr[32706]= 1171527280;
assign addr[32707]= 1106691431;
assign addr[32708]= 1040451659;
assign addr[32709]= 972891995;
assign addr[32710]= 904098143;
assign addr[32711]= 834157373;
assign addr[32712]= 763158411;
assign addr[32713]= 691191324;
assign addr[32714]= 618347408;
assign addr[32715]= 544719071;
assign addr[32716]= 470399716;
assign addr[32717]= 395483624;
assign addr[32718]= 320065829;
assign addr[32719]= 244242007;
assign addr[32720]= 168108346;
assign addr[32721]= 91761426;
assign addr[32722]= 15298099;
assign addr[32723]= -61184634;
assign addr[32724]= -137589750;
assign addr[32725]= -213820322;
assign addr[32726]= -289779648;
assign addr[32727]= -365371365;
assign addr[32728]= -440499581;
assign addr[32729]= -515068990;
assign addr[32730]= -588984994;
assign addr[32731]= -662153826;
assign addr[32732]= -734482665;
assign addr[32733]= -805879757;
assign addr[32734]= -876254528;
assign addr[32735]= -945517704;
assign addr[32736]= -1013581418;
assign addr[32737]= -1080359326;
assign addr[32738]= -1145766716;
assign addr[32739]= -1209720613;
assign addr[32740]= -1272139887;
assign addr[32741]= -1332945355;
assign addr[32742]= -1392059879;
assign addr[32743]= -1449408469;
assign addr[32744]= -1504918373;
assign addr[32745]= -1558519173;
assign addr[32746]= -1610142873;
assign addr[32747]= -1659723983;
assign addr[32748]= -1707199606;
assign addr[32749]= -1752509516;
assign addr[32750]= -1795596234;
assign addr[32751]= -1836405100;
assign addr[32752]= -1874884346;
assign addr[32753]= -1910985158;
assign addr[32754]= -1944661739;
assign addr[32755]= -1975871368;
assign addr[32756]= -2004574453;
assign addr[32757]= -2030734582;
assign addr[32758]= -2054318569;
assign addr[32759]= -2075296495;
assign addr[32760]= -2093641749;
assign addr[32761]= -2109331059;
assign addr[32762]= -2122344521;
assign addr[32763]= -2132665626;
assign addr[32764]= -2140281282;
assign addr[32765]= -2145181827;
assign addr[32766]= -2147361045;
assign addr[32767]= -2146816171;
assign addr[32768]= -2143547897;
assign addr[32769]= -2137560369;
assign addr[32770]= -2128861181;
assign addr[32771]= -2117461370;
assign addr[32772]= -2103375398;
assign addr[32773]= -2086621133;
assign addr[32774]= -2067219829;
assign addr[32775]= -2045196100;
assign addr[32776]= -2020577882;
assign addr[32777]= -1993396407;
assign addr[32778]= -1963686155;
assign addr[32779]= -1931484818;
assign addr[32780]= -1896833245;
assign addr[32781]= -1859775393;
assign addr[32782]= -1820358275;
assign addr[32783]= -1778631892;
assign addr[32784]= -1734649179;
assign addr[32785]= -1688465931;
assign addr[32786]= -1640140734;
assign addr[32787]= -1589734894;
assign addr[32788]= -1537312353;
assign addr[32789]= -1482939614;
assign addr[32790]= -1426685652;
assign addr[32791]= -1368621831;
assign addr[32792]= -1308821808;
assign addr[32793]= -1247361445;
assign addr[32794]= -1184318708;
assign addr[32795]= -1119773573;
assign addr[32796]= -1053807919;
assign addr[32797]= -986505429;
assign addr[32798]= -917951481;
assign addr[32799]= -848233042;
assign addr[32800]= -777438554;
assign addr[32801]= -705657826;
assign addr[32802]= -632981917;
assign addr[32803]= -559503022;
assign addr[32804]= -485314355;
assign addr[32805]= -410510029;
assign addr[32806]= -335184940;
assign addr[32807]= -259434643;
assign addr[32808]= -183355234;
assign addr[32809]= -107043224;
assign addr[32810]= -30595422;
assign addr[32811]= 45891193;
assign addr[32812]= 122319591;
assign addr[32813]= 198592817;
assign addr[32814]= 274614114;
assign addr[32815]= 350287041;
assign addr[32816]= 425515602;
assign addr[32817]= 500204365;
assign addr[32818]= 574258580;
assign addr[32819]= 647584304;
assign addr[32820]= 720088517;
assign addr[32821]= 791679244;
assign addr[32822]= 862265664;
assign addr[32823]= 931758235;
assign addr[32824]= 1000068799;
assign addr[32825]= 1067110699;
assign addr[32826]= 1132798888;
assign addr[32827]= 1197050035;
assign addr[32828]= 1259782632;
assign addr[32829]= 1320917099;
assign addr[32830]= 1380375881;
assign addr[32831]= 1438083551;
assign addr[32832]= 1493966902;
assign addr[32833]= 1547955041;
assign addr[32834]= 1599979481;
assign addr[32835]= 1649974225;
assign addr[32836]= 1697875851;
assign addr[32837]= 1743623590;
assign addr[32838]= 1787159411;
assign addr[32839]= 1828428082;
assign addr[32840]= 1867377253;
assign addr[32841]= 1903957513;
assign addr[32842]= 1938122457;
assign addr[32843]= 1969828744;
assign addr[32844]= 1999036154;
assign addr[32845]= 2025707632;
assign addr[32846]= 2049809346;
assign addr[32847]= 2071310720;
assign addr[32848]= 2090184478;
assign addr[32849]= 2106406677;
assign addr[32850]= 2119956737;
assign addr[32851]= 2130817471;
assign addr[32852]= 2138975100;
assign addr[32853]= 2144419275;
assign addr[32854]= 2147143090;
assign addr[32855]= 2147143090;
assign addr[32856]= 2144419275;
assign addr[32857]= 2138975100;
assign addr[32858]= 2130817471;
assign addr[32859]= 2119956737;
assign addr[32860]= 2106406677;
assign addr[32861]= 2090184478;
assign addr[32862]= 2071310720;
assign addr[32863]= 2049809346;
assign addr[32864]= 2025707632;
assign addr[32865]= 1999036154;
assign addr[32866]= 1969828744;
assign addr[32867]= 1938122457;
assign addr[32868]= 1903957513;
assign addr[32869]= 1867377253;
assign addr[32870]= 1828428082;
assign addr[32871]= 1787159411;
assign addr[32872]= 1743623590;
assign addr[32873]= 1697875851;
assign addr[32874]= 1649974225;
assign addr[32875]= 1599979481;
assign addr[32876]= 1547955041;
assign addr[32877]= 1493966902;
assign addr[32878]= 1438083551;
assign addr[32879]= 1380375881;
assign addr[32880]= 1320917099;
assign addr[32881]= 1259782632;
assign addr[32882]= 1197050035;
assign addr[32883]= 1132798888;
assign addr[32884]= 1067110699;
assign addr[32885]= 1000068799;
assign addr[32886]= 931758235;
assign addr[32887]= 862265664;
assign addr[32888]= 791679244;
assign addr[32889]= 720088517;
assign addr[32890]= 647584304;
assign addr[32891]= 574258580;
assign addr[32892]= 500204365;
assign addr[32893]= 425515602;
assign addr[32894]= 350287041;
assign addr[32895]= 274614114;
assign addr[32896]= 198592817;
assign addr[32897]= 122319591;
assign addr[32898]= 45891193;
assign addr[32899]= -30595422;
assign addr[32900]= -107043224;
assign addr[32901]= -183355234;
assign addr[32902]= -259434643;
assign addr[32903]= -335184940;
assign addr[32904]= -410510029;
assign addr[32905]= -485314355;
assign addr[32906]= -559503022;
assign addr[32907]= -632981917;
assign addr[32908]= -705657826;
assign addr[32909]= -777438554;
assign addr[32910]= -848233042;
assign addr[32911]= -917951481;
assign addr[32912]= -986505429;
assign addr[32913]= -1053807919;
assign addr[32914]= -1119773573;
assign addr[32915]= -1184318708;
assign addr[32916]= -1247361445;
assign addr[32917]= -1308821808;
assign addr[32918]= -1368621831;
assign addr[32919]= -1426685652;
assign addr[32920]= -1482939614;
assign addr[32921]= -1537312353;
assign addr[32922]= -1589734894;
assign addr[32923]= -1640140734;
assign addr[32924]= -1688465931;
assign addr[32925]= -1734649179;
assign addr[32926]= -1778631892;
assign addr[32927]= -1820358275;
assign addr[32928]= -1859775393;
assign addr[32929]= -1896833245;
assign addr[32930]= -1931484818;
assign addr[32931]= -1963686155;
assign addr[32932]= -1993396407;
assign addr[32933]= -2020577882;
assign addr[32934]= -2045196100;
assign addr[32935]= -2067219829;
assign addr[32936]= -2086621133;
assign addr[32937]= -2103375398;
assign addr[32938]= -2117461370;
assign addr[32939]= -2128861181;
assign addr[32940]= -2137560369;
assign addr[32941]= -2143547897;
assign addr[32942]= -2146816171;
assign addr[32943]= -2147361045;
assign addr[32944]= -2145181827;
assign addr[32945]= -2140281282;
assign addr[32946]= -2132665626;
assign addr[32947]= -2122344521;
assign addr[32948]= -2109331059;
assign addr[32949]= -2093641749;
assign addr[32950]= -2075296495;
assign addr[32951]= -2054318569;
assign addr[32952]= -2030734582;
assign addr[32953]= -2004574453;
assign addr[32954]= -1975871368;
assign addr[32955]= -1944661739;
assign addr[32956]= -1910985158;
assign addr[32957]= -1874884346;
assign addr[32958]= -1836405100;
assign addr[32959]= -1795596234;
assign addr[32960]= -1752509516;
assign addr[32961]= -1707199606;
assign addr[32962]= -1659723983;
assign addr[32963]= -1610142873;
assign addr[32964]= -1558519173;
assign addr[32965]= -1504918373;
assign addr[32966]= -1449408469;
assign addr[32967]= -1392059879;
assign addr[32968]= -1332945355;
assign addr[32969]= -1272139887;
assign addr[32970]= -1209720613;
assign addr[32971]= -1145766716;
assign addr[32972]= -1080359326;
assign addr[32973]= -1013581418;
assign addr[32974]= -945517704;
assign addr[32975]= -876254528;
assign addr[32976]= -805879757;
assign addr[32977]= -734482665;
assign addr[32978]= -662153826;
assign addr[32979]= -588984994;
assign addr[32980]= -515068990;
assign addr[32981]= -440499581;
assign addr[32982]= -365371365;
assign addr[32983]= -289779648;
assign addr[32984]= -213820322;
assign addr[32985]= -137589750;
assign addr[32986]= -61184634;
assign addr[32987]= 15298099;
assign addr[32988]= 91761426;
assign addr[32989]= 168108346;
assign addr[32990]= 244242007;
assign addr[32991]= 320065829;
assign addr[32992]= 395483624;
assign addr[32993]= 470399716;
assign addr[32994]= 544719071;
assign addr[32995]= 618347408;
assign addr[32996]= 691191324;
assign addr[32997]= 763158411;
assign addr[32998]= 834157373;
assign addr[32999]= 904098143;
assign addr[33000]= 972891995;
assign addr[33001]= 1040451659;
assign addr[33002]= 1106691431;
assign addr[33003]= 1171527280;
assign addr[33004]= 1234876957;
assign addr[33005]= 1296660098;
assign addr[33006]= 1356798326;
assign addr[33007]= 1415215352;
assign addr[33008]= 1471837070;
assign addr[33009]= 1526591649;
assign addr[33010]= 1579409630;
assign addr[33011]= 1630224009;
assign addr[33012]= 1678970324;
assign addr[33013]= 1725586737;
assign addr[33014]= 1770014111;
assign addr[33015]= 1812196087;
assign addr[33016]= 1852079154;
assign addr[33017]= 1889612716;
assign addr[33018]= 1924749160;
assign addr[33019]= 1957443913;
assign addr[33020]= 1987655498;
assign addr[33021]= 2015345591;
assign addr[33022]= 2040479063;
assign addr[33023]= 2063024031;
assign addr[33024]= 2082951896;
assign addr[33025]= 2100237377;
assign addr[33026]= 2114858546;
assign addr[33027]= 2126796855;
assign addr[33028]= 2136037160;
assign addr[33029]= 2142567738;
assign addr[33030]= 2146380306;
assign addr[33031]= 2147470025;
assign addr[33032]= 2145835515;
assign addr[33033]= 2141478848;
assign addr[33034]= 2134405552;
assign addr[33035]= 2124624598;
assign addr[33036]= 2112148396;
assign addr[33037]= 2096992772;
assign addr[33038]= 2079176953;
assign addr[33039]= 2058723538;
assign addr[33040]= 2035658475;
assign addr[33041]= 2010011024;
assign addr[33042]= 1981813720;
assign addr[33043]= 1951102334;
assign addr[33044]= 1917915825;
assign addr[33045]= 1882296293;
assign addr[33046]= 1844288924;
assign addr[33047]= 1803941934;
assign addr[33048]= 1761306505;
assign addr[33049]= 1716436725;
assign addr[33050]= 1669389513;
assign addr[33051]= 1620224553;
assign addr[33052]= 1569004214;
assign addr[33053]= 1515793473;
assign addr[33054]= 1460659832;
assign addr[33055]= 1403673233;
assign addr[33056]= 1344905966;
assign addr[33057]= 1284432584;
assign addr[33058]= 1222329801;
assign addr[33059]= 1158676398;
assign addr[33060]= 1093553126;
assign addr[33061]= 1027042599;
assign addr[33062]= 959229189;
assign addr[33063]= 890198924;
assign addr[33064]= 820039373;
assign addr[33065]= 748839539;
assign addr[33066]= 676689746;
assign addr[33067]= 603681519;
assign addr[33068]= 529907477;
assign addr[33069]= 455461206;
assign addr[33070]= 380437148;
assign addr[33071]= 304930476;
assign addr[33072]= 229036977;
assign addr[33073]= 152852926;
assign addr[33074]= 76474970;
assign addr[33075]= 0;
assign addr[33076]= -76474970;
assign addr[33077]= -152852926;
assign addr[33078]= -229036977;
assign addr[33079]= -304930476;
assign addr[33080]= -380437148;
assign addr[33081]= -455461206;
assign addr[33082]= -529907477;
assign addr[33083]= -603681519;
assign addr[33084]= -676689746;
assign addr[33085]= -748839539;
assign addr[33086]= -820039373;
assign addr[33087]= -890198924;
assign addr[33088]= -959229189;
assign addr[33089]= -1027042599;
assign addr[33090]= -1093553126;
assign addr[33091]= -1158676398;
assign addr[33092]= -1222329801;
assign addr[33093]= -1284432584;
assign addr[33094]= -1344905966;
assign addr[33095]= -1403673233;
assign addr[33096]= -1460659832;
assign addr[33097]= -1515793473;
assign addr[33098]= -1569004214;
assign addr[33099]= -1620224553;
assign addr[33100]= -1669389513;
assign addr[33101]= -1716436725;
assign addr[33102]= -1761306505;
assign addr[33103]= -1803941934;
assign addr[33104]= -1844288924;
assign addr[33105]= -1882296293;
assign addr[33106]= -1917915825;
assign addr[33107]= -1951102334;
assign addr[33108]= -1981813720;
assign addr[33109]= -2010011024;
assign addr[33110]= -2035658475;
assign addr[33111]= -2058723538;
assign addr[33112]= -2079176953;
assign addr[33113]= -2096992772;
assign addr[33114]= -2112148396;
assign addr[33115]= -2124624598;
assign addr[33116]= -2134405552;
assign addr[33117]= -2141478848;
assign addr[33118]= -2145835515;
assign addr[33119]= -2147470025;
assign addr[33120]= -2146380306;
assign addr[33121]= -2142567738;
assign addr[33122]= -2136037160;
assign addr[33123]= -2126796855;
assign addr[33124]= -2114858546;
assign addr[33125]= -2100237377;
assign addr[33126]= -2082951896;
assign addr[33127]= -2063024031;
assign addr[33128]= -2040479063;
assign addr[33129]= -2015345591;
assign addr[33130]= -1987655498;
assign addr[33131]= -1957443913;
assign addr[33132]= -1924749160;
assign addr[33133]= -1889612716;
assign addr[33134]= -1852079154;
assign addr[33135]= -1812196087;
assign addr[33136]= -1770014111;
assign addr[33137]= -1725586737;
assign addr[33138]= -1678970324;
assign addr[33139]= -1630224009;
assign addr[33140]= -1579409630;
assign addr[33141]= -1526591649;
assign addr[33142]= -1471837070;
assign addr[33143]= -1415215352;
assign addr[33144]= -1356798326;
assign addr[33145]= -1296660098;
assign addr[33146]= -1234876957;
assign addr[33147]= -1171527280;
assign addr[33148]= -1106691431;
assign addr[33149]= -1040451659;
assign addr[33150]= -972891995;
assign addr[33151]= -904098143;
assign addr[33152]= -834157373;
assign addr[33153]= -763158411;
assign addr[33154]= -691191324;
assign addr[33155]= -618347408;
assign addr[33156]= -544719071;
assign addr[33157]= -470399716;
assign addr[33158]= -395483624;
assign addr[33159]= -320065829;
assign addr[33160]= -244242007;
assign addr[33161]= -168108346;
assign addr[33162]= -91761426;
assign addr[33163]= -15298099;
assign addr[33164]= 61184634;
assign addr[33165]= 137589750;
assign addr[33166]= 213820322;
assign addr[33167]= 289779648;
assign addr[33168]= 365371365;
assign addr[33169]= 440499581;
assign addr[33170]= 515068990;
assign addr[33171]= 588984994;
assign addr[33172]= 662153826;
assign addr[33173]= 734482665;
assign addr[33174]= 805879757;
assign addr[33175]= 876254528;
assign addr[33176]= 945517704;
assign addr[33177]= 1013581418;
assign addr[33178]= 1080359326;
assign addr[33179]= 1145766716;
assign addr[33180]= 1209720613;
assign addr[33181]= 1272139887;
assign addr[33182]= 1332945355;
assign addr[33183]= 1392059879;
assign addr[33184]= 1449408469;
assign addr[33185]= 1504918373;
assign addr[33186]= 1558519173;
assign addr[33187]= 1610142873;
assign addr[33188]= 1659723983;
assign addr[33189]= 1707199606;
assign addr[33190]= 1752509516;
assign addr[33191]= 1795596234;
assign addr[33192]= 1836405100;
assign addr[33193]= 1874884346;
assign addr[33194]= 1910985158;
assign addr[33195]= 1944661739;
assign addr[33196]= 1975871368;
assign addr[33197]= 2004574453;
assign addr[33198]= 2030734582;
assign addr[33199]= 2054318569;
assign addr[33200]= 2075296495;
assign addr[33201]= 2093641749;
assign addr[33202]= 2109331059;
assign addr[33203]= 2122344521;
assign addr[33204]= 2132665626;
assign addr[33205]= 2140281282;
assign addr[33206]= 2145181827;
assign addr[33207]= 2147361045;
assign addr[33208]= 2146816171;
assign addr[33209]= 2143547897;
assign addr[33210]= 2137560369;
assign addr[33211]= 2128861181;
assign addr[33212]= 2117461370;
assign addr[33213]= 2103375398;
assign addr[33214]= 2086621133;
assign addr[33215]= 2067219829;
assign addr[33216]= 2045196100;
assign addr[33217]= 2020577882;
assign addr[33218]= 1993396407;
assign addr[33219]= 1963686155;
assign addr[33220]= 1931484818;
assign addr[33221]= 1896833245;
assign addr[33222]= 1859775393;
assign addr[33223]= 1820358275;
assign addr[33224]= 1778631892;
assign addr[33225]= 1734649179;
assign addr[33226]= 1688465931;
assign addr[33227]= 1640140734;
assign addr[33228]= 1589734894;
assign addr[33229]= 1537312353;
assign addr[33230]= 1482939614;
assign addr[33231]= 1426685652;
assign addr[33232]= 1368621831;
assign addr[33233]= 1308821808;
assign addr[33234]= 1247361445;
assign addr[33235]= 1184318708;
assign addr[33236]= 1119773573;
assign addr[33237]= 1053807919;
assign addr[33238]= 986505429;
assign addr[33239]= 917951481;
assign addr[33240]= 848233042;
assign addr[33241]= 777438554;
assign addr[33242]= 705657826;
assign addr[33243]= 632981917;
assign addr[33244]= 559503022;
assign addr[33245]= 485314355;
assign addr[33246]= 410510029;
assign addr[33247]= 335184940;
assign addr[33248]= 259434643;
assign addr[33249]= 183355234;
assign addr[33250]= 107043224;
assign addr[33251]= 30595422;
assign addr[33252]= -45891193;
assign addr[33253]= -122319591;
assign addr[33254]= -198592817;
assign addr[33255]= -274614114;
assign addr[33256]= -350287041;
assign addr[33257]= -425515602;
assign addr[33258]= -500204365;
assign addr[33259]= -574258580;
assign addr[33260]= -647584304;
assign addr[33261]= -720088517;
assign addr[33262]= -791679244;
assign addr[33263]= -862265664;
assign addr[33264]= -931758235;
assign addr[33265]= -1000068799;
assign addr[33266]= -1067110699;
assign addr[33267]= -1132798888;
assign addr[33268]= -1197050035;
assign addr[33269]= -1259782632;
assign addr[33270]= -1320917099;
assign addr[33271]= -1380375881;
assign addr[33272]= -1438083551;
assign addr[33273]= -1493966902;
assign addr[33274]= -1547955041;
assign addr[33275]= -1599979481;
assign addr[33276]= -1649974225;
assign addr[33277]= -1697875851;
assign addr[33278]= -1743623590;
assign addr[33279]= -1787159411;
assign addr[33280]= -1828428082;
assign addr[33281]= -1867377253;
assign addr[33282]= -1903957513;
assign addr[33283]= -1938122457;
assign addr[33284]= -1969828744;
assign addr[33285]= -1999036154;
assign addr[33286]= -2025707632;
assign addr[33287]= -2049809346;
assign addr[33288]= -2071310720;
assign addr[33289]= -2090184478;
assign addr[33290]= -2106406677;
assign addr[33291]= -2119956737;
assign addr[33292]= -2130817471;
assign addr[33293]= -2138975100;
assign addr[33294]= -2144419275;
assign addr[33295]= -2147143090;
assign addr[33296]= -2147143090;
assign addr[33297]= -2144419275;
assign addr[33298]= -2138975100;
assign addr[33299]= -2130817471;
assign addr[33300]= -2119956737;
assign addr[33301]= -2106406677;
assign addr[33302]= -2090184478;
assign addr[33303]= -2071310720;
assign addr[33304]= -2049809346;
assign addr[33305]= -2025707632;
assign addr[33306]= -1999036154;
assign addr[33307]= -1969828744;
assign addr[33308]= -1938122457;
assign addr[33309]= -1903957513;
assign addr[33310]= -1867377253;
assign addr[33311]= -1828428082;
assign addr[33312]= -1787159411;
assign addr[33313]= -1743623590;
assign addr[33314]= -1697875851;
assign addr[33315]= -1649974225;
assign addr[33316]= -1599979481;
assign addr[33317]= -1547955041;
assign addr[33318]= -1493966902;
assign addr[33319]= -1438083551;
assign addr[33320]= -1380375881;
assign addr[33321]= -1320917099;
assign addr[33322]= -1259782632;
assign addr[33323]= -1197050035;
assign addr[33324]= -1132798888;
assign addr[33325]= -1067110699;
assign addr[33326]= -1000068799;
assign addr[33327]= -931758235;
assign addr[33328]= -862265664;
assign addr[33329]= -791679244;
assign addr[33330]= -720088517;
assign addr[33331]= -647584304;
assign addr[33332]= -574258580;
assign addr[33333]= -500204365;
assign addr[33334]= -425515602;
assign addr[33335]= -350287041;
assign addr[33336]= -274614114;
assign addr[33337]= -198592817;
assign addr[33338]= -122319591;
assign addr[33339]= -45891193;
assign addr[33340]= 30595422;
assign addr[33341]= 107043224;
assign addr[33342]= 183355234;
assign addr[33343]= 259434643;
assign addr[33344]= 335184940;
assign addr[33345]= 410510029;
assign addr[33346]= 485314355;
assign addr[33347]= 559503022;
assign addr[33348]= 632981917;
assign addr[33349]= 705657826;
assign addr[33350]= 777438554;
assign addr[33351]= 848233042;
assign addr[33352]= 917951481;
assign addr[33353]= 986505429;
assign addr[33354]= 1053807919;
assign addr[33355]= 1119773573;
assign addr[33356]= 1184318708;
assign addr[33357]= 1247361445;
assign addr[33358]= 1308821808;
assign addr[33359]= 1368621831;
assign addr[33360]= 1426685652;
assign addr[33361]= 1482939614;
assign addr[33362]= 1537312353;
assign addr[33363]= 1589734894;
assign addr[33364]= 1640140734;
assign addr[33365]= 1688465931;
assign addr[33366]= 1734649179;
assign addr[33367]= 1778631892;
assign addr[33368]= 1820358275;
assign addr[33369]= 1859775393;
assign addr[33370]= 1896833245;
assign addr[33371]= 1931484818;
assign addr[33372]= 1963686155;
assign addr[33373]= 1993396407;
assign addr[33374]= 2020577882;
assign addr[33375]= 2045196100;
assign addr[33376]= 2067219829;
assign addr[33377]= 2086621133;
assign addr[33378]= 2103375398;
assign addr[33379]= 2117461370;
assign addr[33380]= 2128861181;
assign addr[33381]= 2137560369;
assign addr[33382]= 2143547897;
assign addr[33383]= 2146816171;
assign addr[33384]= 2147361045;
assign addr[33385]= 2145181827;
assign addr[33386]= 2140281282;
assign addr[33387]= 2132665626;
assign addr[33388]= 2122344521;
assign addr[33389]= 2109331059;
assign addr[33390]= 2093641749;
assign addr[33391]= 2075296495;
assign addr[33392]= 2054318569;
assign addr[33393]= 2030734582;
assign addr[33394]= 2004574453;
assign addr[33395]= 1975871368;
assign addr[33396]= 1944661739;
assign addr[33397]= 1910985158;
assign addr[33398]= 1874884346;
assign addr[33399]= 1836405100;
assign addr[33400]= 1795596234;
assign addr[33401]= 1752509516;
assign addr[33402]= 1707199606;
assign addr[33403]= 1659723983;
assign addr[33404]= 1610142873;
assign addr[33405]= 1558519173;
assign addr[33406]= 1504918373;
assign addr[33407]= 1449408469;
assign addr[33408]= 1392059879;
assign addr[33409]= 1332945355;
assign addr[33410]= 1272139887;
assign addr[33411]= 1209720613;
assign addr[33412]= 1145766716;
assign addr[33413]= 1080359326;
assign addr[33414]= 1013581418;
assign addr[33415]= 945517704;
assign addr[33416]= 876254528;
assign addr[33417]= 805879757;
assign addr[33418]= 734482665;
assign addr[33419]= 662153826;
assign addr[33420]= 588984994;
assign addr[33421]= 515068990;
assign addr[33422]= 440499581;
assign addr[33423]= 365371365;
assign addr[33424]= 289779648;
assign addr[33425]= 213820322;
assign addr[33426]= 137589750;
assign addr[33427]= 61184634;
assign addr[33428]= -15298099;
assign addr[33429]= -91761426;
assign addr[33430]= -168108346;
assign addr[33431]= -244242007;
assign addr[33432]= -320065829;
assign addr[33433]= -395483624;
assign addr[33434]= -470399716;
assign addr[33435]= -544719071;
assign addr[33436]= -618347408;
assign addr[33437]= -691191324;
assign addr[33438]= -763158411;
assign addr[33439]= -834157373;
assign addr[33440]= -904098143;
assign addr[33441]= -972891995;
assign addr[33442]= -1040451659;
assign addr[33443]= -1106691431;
assign addr[33444]= -1171527280;
assign addr[33445]= -1234876957;
assign addr[33446]= -1296660098;
assign addr[33447]= -1356798326;
assign addr[33448]= -1415215352;
assign addr[33449]= -1471837070;
assign addr[33450]= -1526591649;
assign addr[33451]= -1579409630;
assign addr[33452]= -1630224009;
assign addr[33453]= -1678970324;
assign addr[33454]= -1725586737;
assign addr[33455]= -1770014111;
assign addr[33456]= -1812196087;
assign addr[33457]= -1852079154;
assign addr[33458]= -1889612716;
assign addr[33459]= -1924749160;
assign addr[33460]= -1957443913;
assign addr[33461]= -1987655498;
assign addr[33462]= -2015345591;
assign addr[33463]= -2040479063;
assign addr[33464]= -2063024031;
assign addr[33465]= -2082951896;
assign addr[33466]= -2100237377;
assign addr[33467]= -2114858546;
assign addr[33468]= -2126796855;
assign addr[33469]= -2136037160;
assign addr[33470]= -2142567738;
assign addr[33471]= -2146380306;
assign addr[33472]= -2147470025;
assign addr[33473]= -2145835515;
assign addr[33474]= -2141478848;
assign addr[33475]= -2134405552;
assign addr[33476]= -2124624598;
assign addr[33477]= -2112148396;
assign addr[33478]= -2096992772;
assign addr[33479]= -2079176953;
assign addr[33480]= -2058723538;
assign addr[33481]= -2035658475;
assign addr[33482]= -2010011024;
assign addr[33483]= -1981813720;
assign addr[33484]= -1951102334;
assign addr[33485]= -1917915825;
assign addr[33486]= -1882296293;
assign addr[33487]= -1844288924;
assign addr[33488]= -1803941934;
assign addr[33489]= -1761306505;
assign addr[33490]= -1716436725;
assign addr[33491]= -1669389513;
assign addr[33492]= -1620224553;
assign addr[33493]= -1569004214;
assign addr[33494]= -1515793473;
assign addr[33495]= -1460659832;
assign addr[33496]= -1403673233;
assign addr[33497]= -1344905966;
assign addr[33498]= -1284432584;
assign addr[33499]= -1222329801;
assign addr[33500]= -1158676398;
assign addr[33501]= -1093553126;
assign addr[33502]= -1027042599;
assign addr[33503]= -959229189;
assign addr[33504]= -890198924;
assign addr[33505]= -820039373;
assign addr[33506]= -748839539;
assign addr[33507]= -676689746;
assign addr[33508]= -603681519;
assign addr[33509]= -529907477;
assign addr[33510]= -455461206;
assign addr[33511]= -380437148;
assign addr[33512]= -304930476;
assign addr[33513]= -229036977;
assign addr[33514]= -152852926;
assign addr[33515]= -76474970;
assign addr[33516]= 0;
assign addr[33517]= 76474970;
assign addr[33518]= 152852926;
assign addr[33519]= 229036977;
assign addr[33520]= 304930476;
assign addr[33521]= 380437148;
assign addr[33522]= 455461206;
assign addr[33523]= 529907477;
assign addr[33524]= 603681519;
assign addr[33525]= 676689746;
assign addr[33526]= 748839539;
assign addr[33527]= 820039373;
assign addr[33528]= 890198924;
assign addr[33529]= 959229189;
assign addr[33530]= 1027042599;
assign addr[33531]= 1093553126;
assign addr[33532]= 1158676398;
assign addr[33533]= 1222329801;
assign addr[33534]= 1284432584;
assign addr[33535]= 1344905966;
assign addr[33536]= 1403673233;
assign addr[33537]= 1460659832;
assign addr[33538]= 1515793473;
assign addr[33539]= 1569004214;
assign addr[33540]= 1620224553;
assign addr[33541]= 1669389513;
assign addr[33542]= 1716436725;
assign addr[33543]= 1761306505;
assign addr[33544]= 1803941934;
assign addr[33545]= 1844288924;
assign addr[33546]= 1882296293;
assign addr[33547]= 1917915825;
assign addr[33548]= 1951102334;
assign addr[33549]= 1981813720;
assign addr[33550]= 2010011024;
assign addr[33551]= 2035658475;
assign addr[33552]= 2058723538;
assign addr[33553]= 2079176953;
assign addr[33554]= 2096992772;
assign addr[33555]= 2112148396;
assign addr[33556]= 2124624598;
assign addr[33557]= 2134405552;
assign addr[33558]= 2141478848;
assign addr[33559]= 2145835515;
assign addr[33560]= 2147470025;
assign addr[33561]= 2146380306;
assign addr[33562]= 2142567738;
assign addr[33563]= 2136037160;
assign addr[33564]= 2126796855;
assign addr[33565]= 2114858546;
assign addr[33566]= 2100237377;
assign addr[33567]= 2082951896;
assign addr[33568]= 2063024031;
assign addr[33569]= 2040479063;
assign addr[33570]= 2015345591;
assign addr[33571]= 1987655498;
assign addr[33572]= 1957443913;
assign addr[33573]= 1924749160;
assign addr[33574]= 1889612716;
assign addr[33575]= 1852079154;
assign addr[33576]= 1812196087;
assign addr[33577]= 1770014111;
assign addr[33578]= 1725586737;
assign addr[33579]= 1678970324;
assign addr[33580]= 1630224009;
assign addr[33581]= 1579409630;
assign addr[33582]= 1526591649;
assign addr[33583]= 1471837070;
assign addr[33584]= 1415215352;
assign addr[33585]= 1356798326;
assign addr[33586]= 1296660098;
assign addr[33587]= 1234876957;
assign addr[33588]= 1171527280;
assign addr[33589]= 1106691431;
assign addr[33590]= 1040451659;
assign addr[33591]= 972891995;
assign addr[33592]= 904098143;
assign addr[33593]= 834157373;
assign addr[33594]= 763158411;
assign addr[33595]= 691191324;
assign addr[33596]= 618347408;
assign addr[33597]= 544719071;
assign addr[33598]= 470399716;
assign addr[33599]= 395483624;
assign addr[33600]= 320065829;
assign addr[33601]= 244242007;
assign addr[33602]= 168108346;
assign addr[33603]= 91761426;
assign addr[33604]= 15298099;
assign addr[33605]= -61184634;
assign addr[33606]= -137589750;
assign addr[33607]= -213820322;
assign addr[33608]= -289779648;
assign addr[33609]= -365371365;
assign addr[33610]= -440499581;
assign addr[33611]= -515068990;
assign addr[33612]= -588984994;
assign addr[33613]= -662153826;
assign addr[33614]= -734482665;
assign addr[33615]= -805879757;
assign addr[33616]= -876254528;
assign addr[33617]= -945517704;
assign addr[33618]= -1013581418;
assign addr[33619]= -1080359326;
assign addr[33620]= -1145766716;
assign addr[33621]= -1209720613;
assign addr[33622]= -1272139887;
assign addr[33623]= -1332945355;
assign addr[33624]= -1392059879;
assign addr[33625]= -1449408469;
assign addr[33626]= -1504918373;
assign addr[33627]= -1558519173;
assign addr[33628]= -1610142873;
assign addr[33629]= -1659723983;
assign addr[33630]= -1707199606;
assign addr[33631]= -1752509516;
assign addr[33632]= -1795596234;
assign addr[33633]= -1836405100;
assign addr[33634]= -1874884346;
assign addr[33635]= -1910985158;
assign addr[33636]= -1944661739;
assign addr[33637]= -1975871368;
assign addr[33638]= -2004574453;
assign addr[33639]= -2030734582;
assign addr[33640]= -2054318569;
assign addr[33641]= -2075296495;
assign addr[33642]= -2093641749;
assign addr[33643]= -2109331059;
assign addr[33644]= -2122344521;
assign addr[33645]= -2132665626;
assign addr[33646]= -2140281282;
assign addr[33647]= -2145181827;
assign addr[33648]= -2147361045;
assign addr[33649]= -2146816171;
assign addr[33650]= -2143547897;
assign addr[33651]= -2137560369;
assign addr[33652]= -2128861181;
assign addr[33653]= -2117461370;
assign addr[33654]= -2103375398;
assign addr[33655]= -2086621133;
assign addr[33656]= -2067219829;
assign addr[33657]= -2045196100;
assign addr[33658]= -2020577882;
assign addr[33659]= -1993396407;
assign addr[33660]= -1963686155;
assign addr[33661]= -1931484818;
assign addr[33662]= -1896833245;
assign addr[33663]= -1859775393;
assign addr[33664]= -1820358275;
assign addr[33665]= -1778631892;
assign addr[33666]= -1734649179;
assign addr[33667]= -1688465931;
assign addr[33668]= -1640140734;
assign addr[33669]= -1589734894;
assign addr[33670]= -1537312353;
assign addr[33671]= -1482939614;
assign addr[33672]= -1426685652;
assign addr[33673]= -1368621831;
assign addr[33674]= -1308821808;
assign addr[33675]= -1247361445;
assign addr[33676]= -1184318708;
assign addr[33677]= -1119773573;
assign addr[33678]= -1053807919;
assign addr[33679]= -986505429;
assign addr[33680]= -917951481;
assign addr[33681]= -848233042;
assign addr[33682]= -777438554;
assign addr[33683]= -705657826;
assign addr[33684]= -632981917;
assign addr[33685]= -559503022;
assign addr[33686]= -485314355;
assign addr[33687]= -410510029;
assign addr[33688]= -335184940;
assign addr[33689]= -259434643;
assign addr[33690]= -183355234;
assign addr[33691]= -107043224;
assign addr[33692]= -30595422;
assign addr[33693]= 45891193;
assign addr[33694]= 122319591;
assign addr[33695]= 198592817;
assign addr[33696]= 274614114;
assign addr[33697]= 350287041;
assign addr[33698]= 425515602;
assign addr[33699]= 500204365;
assign addr[33700]= 574258580;
assign addr[33701]= 647584304;
assign addr[33702]= 720088517;
assign addr[33703]= 791679244;
assign addr[33704]= 862265664;
assign addr[33705]= 931758235;
assign addr[33706]= 1000068799;
assign addr[33707]= 1067110699;
assign addr[33708]= 1132798888;
assign addr[33709]= 1197050035;
assign addr[33710]= 1259782632;
assign addr[33711]= 1320917099;
assign addr[33712]= 1380375881;
assign addr[33713]= 1438083551;
assign addr[33714]= 1493966902;
assign addr[33715]= 1547955041;
assign addr[33716]= 1599979481;
assign addr[33717]= 1649974225;
assign addr[33718]= 1697875851;
assign addr[33719]= 1743623590;
assign addr[33720]= 1787159411;
assign addr[33721]= 1828428082;
assign addr[33722]= 1867377253;
assign addr[33723]= 1903957513;
assign addr[33724]= 1938122457;
assign addr[33725]= 1969828744;
assign addr[33726]= 1999036154;
assign addr[33727]= 2025707632;
assign addr[33728]= 2049809346;
assign addr[33729]= 2071310720;
assign addr[33730]= 2090184478;
assign addr[33731]= 2106406677;
assign addr[33732]= 2119956737;
assign addr[33733]= 2130817471;
assign addr[33734]= 2138975100;
assign addr[33735]= 2144419275;
assign addr[33736]= 2147143090;
assign addr[33737]= 2147143090;
assign addr[33738]= 2144419275;
assign addr[33739]= 2138975100;
assign addr[33740]= 2130817471;
assign addr[33741]= 2119956737;
assign addr[33742]= 2106406677;
assign addr[33743]= 2090184478;
assign addr[33744]= 2071310720;
assign addr[33745]= 2049809346;
assign addr[33746]= 2025707632;
assign addr[33747]= 1999036154;
assign addr[33748]= 1969828744;
assign addr[33749]= 1938122457;
assign addr[33750]= 1903957513;
assign addr[33751]= 1867377253;
assign addr[33752]= 1828428082;
assign addr[33753]= 1787159411;
assign addr[33754]= 1743623590;
assign addr[33755]= 1697875851;
assign addr[33756]= 1649974225;
assign addr[33757]= 1599979481;
assign addr[33758]= 1547955041;
assign addr[33759]= 1493966902;
assign addr[33760]= 1438083551;
assign addr[33761]= 1380375881;
assign addr[33762]= 1320917099;
assign addr[33763]= 1259782632;
assign addr[33764]= 1197050035;
assign addr[33765]= 1132798888;
assign addr[33766]= 1067110699;
assign addr[33767]= 1000068799;
assign addr[33768]= 931758235;
assign addr[33769]= 862265664;
assign addr[33770]= 791679244;
assign addr[33771]= 720088517;
assign addr[33772]= 647584304;
assign addr[33773]= 574258580;
assign addr[33774]= 500204365;
assign addr[33775]= 425515602;
assign addr[33776]= 350287041;
assign addr[33777]= 274614114;
assign addr[33778]= 198592817;
assign addr[33779]= 122319591;
assign addr[33780]= 45891193;
assign addr[33781]= -30595422;
assign addr[33782]= -107043224;
assign addr[33783]= -183355234;
assign addr[33784]= -259434643;
assign addr[33785]= -335184940;
assign addr[33786]= -410510029;
assign addr[33787]= -485314355;
assign addr[33788]= -559503022;
assign addr[33789]= -632981917;
assign addr[33790]= -705657826;
assign addr[33791]= -777438554;
assign addr[33792]= -848233042;
assign addr[33793]= -917951481;
assign addr[33794]= -986505429;
assign addr[33795]= -1053807919;
assign addr[33796]= -1119773573;
assign addr[33797]= -1184318708;
assign addr[33798]= -1247361445;
assign addr[33799]= -1308821808;
assign addr[33800]= -1368621831;
assign addr[33801]= -1426685652;
assign addr[33802]= -1482939614;
assign addr[33803]= -1537312353;
assign addr[33804]= -1589734894;
assign addr[33805]= -1640140734;
assign addr[33806]= -1688465931;
assign addr[33807]= -1734649179;
assign addr[33808]= -1778631892;
assign addr[33809]= -1820358275;
assign addr[33810]= -1859775393;
assign addr[33811]= -1896833245;
assign addr[33812]= -1931484818;
assign addr[33813]= -1963686155;
assign addr[33814]= -1993396407;
assign addr[33815]= -2020577882;
assign addr[33816]= -2045196100;
assign addr[33817]= -2067219829;
assign addr[33818]= -2086621133;
assign addr[33819]= -2103375398;
assign addr[33820]= -2117461370;
assign addr[33821]= -2128861181;
assign addr[33822]= -2137560369;
assign addr[33823]= -2143547897;
assign addr[33824]= -2146816171;
assign addr[33825]= -2147361045;
assign addr[33826]= -2145181827;
assign addr[33827]= -2140281282;
assign addr[33828]= -2132665626;
assign addr[33829]= -2122344521;
assign addr[33830]= -2109331059;
assign addr[33831]= -2093641749;
assign addr[33832]= -2075296495;
assign addr[33833]= -2054318569;
assign addr[33834]= -2030734582;
assign addr[33835]= -2004574453;
assign addr[33836]= -1975871368;
assign addr[33837]= -1944661739;
assign addr[33838]= -1910985158;
assign addr[33839]= -1874884346;
assign addr[33840]= -1836405100;
assign addr[33841]= -1795596234;
assign addr[33842]= -1752509516;
assign addr[33843]= -1707199606;
assign addr[33844]= -1659723983;
assign addr[33845]= -1610142873;
assign addr[33846]= -1558519173;
assign addr[33847]= -1504918373;
assign addr[33848]= -1449408469;
assign addr[33849]= -1392059879;
assign addr[33850]= -1332945355;
assign addr[33851]= -1272139887;
assign addr[33852]= -1209720613;
assign addr[33853]= -1145766716;
assign addr[33854]= -1080359326;
assign addr[33855]= -1013581418;
assign addr[33856]= -945517704;
assign addr[33857]= -876254528;
assign addr[33858]= -805879757;
assign addr[33859]= -734482665;
assign addr[33860]= -662153826;
assign addr[33861]= -588984994;
assign addr[33862]= -515068990;
assign addr[33863]= -440499581;
assign addr[33864]= -365371365;
assign addr[33865]= -289779648;
assign addr[33866]= -213820322;
assign addr[33867]= -137589750;
assign addr[33868]= -61184634;
assign addr[33869]= 15298099;
assign addr[33870]= 91761426;
assign addr[33871]= 168108346;
assign addr[33872]= 244242007;
assign addr[33873]= 320065829;
assign addr[33874]= 395483624;
assign addr[33875]= 470399716;
assign addr[33876]= 544719071;
assign addr[33877]= 618347408;
assign addr[33878]= 691191324;
assign addr[33879]= 763158411;
assign addr[33880]= 834157373;
assign addr[33881]= 904098143;
assign addr[33882]= 972891995;
assign addr[33883]= 1040451659;
assign addr[33884]= 1106691431;
assign addr[33885]= 1171527280;
assign addr[33886]= 1234876957;
assign addr[33887]= 1296660098;
assign addr[33888]= 1356798326;
assign addr[33889]= 1415215352;
assign addr[33890]= 1471837070;
assign addr[33891]= 1526591649;
assign addr[33892]= 1579409630;
assign addr[33893]= 1630224009;
assign addr[33894]= 1678970324;
assign addr[33895]= 1725586737;
assign addr[33896]= 1770014111;
assign addr[33897]= 1812196087;
assign addr[33898]= 1852079154;
assign addr[33899]= 1889612716;
assign addr[33900]= 1924749160;
assign addr[33901]= 1957443913;
assign addr[33902]= 1987655498;
assign addr[33903]= 2015345591;
assign addr[33904]= 2040479063;
assign addr[33905]= 2063024031;
assign addr[33906]= 2082951896;
assign addr[33907]= 2100237377;
assign addr[33908]= 2114858546;
assign addr[33909]= 2126796855;
assign addr[33910]= 2136037160;
assign addr[33911]= 2142567738;
assign addr[33912]= 2146380306;
assign addr[33913]= 2147470025;
assign addr[33914]= 2145835515;
assign addr[33915]= 2141478848;
assign addr[33916]= 2134405552;
assign addr[33917]= 2124624598;
assign addr[33918]= 2112148396;
assign addr[33919]= 2096992772;
assign addr[33920]= 2079176953;
assign addr[33921]= 2058723538;
assign addr[33922]= 2035658475;
assign addr[33923]= 2010011024;
assign addr[33924]= 1981813720;
assign addr[33925]= 1951102334;
assign addr[33926]= 1917915825;
assign addr[33927]= 1882296293;
assign addr[33928]= 1844288924;
assign addr[33929]= 1803941934;
assign addr[33930]= 1761306505;
assign addr[33931]= 1716436725;
assign addr[33932]= 1669389513;
assign addr[33933]= 1620224553;
assign addr[33934]= 1569004214;
assign addr[33935]= 1515793473;
assign addr[33936]= 1460659832;
assign addr[33937]= 1403673233;
assign addr[33938]= 1344905966;
assign addr[33939]= 1284432584;
assign addr[33940]= 1222329801;
assign addr[33941]= 1158676398;
assign addr[33942]= 1093553126;
assign addr[33943]= 1027042599;
assign addr[33944]= 959229189;
assign addr[33945]= 890198924;
assign addr[33946]= 820039373;
assign addr[33947]= 748839539;
assign addr[33948]= 676689746;
assign addr[33949]= 603681519;
assign addr[33950]= 529907477;
assign addr[33951]= 455461206;
assign addr[33952]= 380437148;
assign addr[33953]= 304930476;
assign addr[33954]= 229036977;
assign addr[33955]= 152852926;
assign addr[33956]= 76474970;
assign addr[33957]= 0;
assign addr[33958]= -76474970;
assign addr[33959]= -152852926;
assign addr[33960]= -229036977;
assign addr[33961]= -304930476;
assign addr[33962]= -380437148;
assign addr[33963]= -455461206;
assign addr[33964]= -529907477;
assign addr[33965]= -603681519;
assign addr[33966]= -676689746;
assign addr[33967]= -748839539;
assign addr[33968]= -820039373;
assign addr[33969]= -890198924;
assign addr[33970]= -959229189;
assign addr[33971]= -1027042599;
assign addr[33972]= -1093553126;
assign addr[33973]= -1158676398;
assign addr[33974]= -1222329801;
assign addr[33975]= -1284432584;
assign addr[33976]= -1344905966;
assign addr[33977]= -1403673233;
assign addr[33978]= -1460659832;
assign addr[33979]= -1515793473;
assign addr[33980]= -1569004214;
assign addr[33981]= -1620224553;
assign addr[33982]= -1669389513;
assign addr[33983]= -1716436725;
assign addr[33984]= -1761306505;
assign addr[33985]= -1803941934;
assign addr[33986]= -1844288924;
assign addr[33987]= -1882296293;
assign addr[33988]= -1917915825;
assign addr[33989]= -1951102334;
assign addr[33990]= -1981813720;
assign addr[33991]= -2010011024;
assign addr[33992]= -2035658475;
assign addr[33993]= -2058723538;
assign addr[33994]= -2079176953;
assign addr[33995]= -2096992772;
assign addr[33996]= -2112148396;
assign addr[33997]= -2124624598;
assign addr[33998]= -2134405552;
assign addr[33999]= -2141478848;
assign addr[34000]= -2145835515;
assign addr[34001]= -2147470025;
assign addr[34002]= -2146380306;
assign addr[34003]= -2142567738;
assign addr[34004]= -2136037160;
assign addr[34005]= -2126796855;
assign addr[34006]= -2114858546;
assign addr[34007]= -2100237377;
assign addr[34008]= -2082951896;
assign addr[34009]= -2063024031;
assign addr[34010]= -2040479063;
assign addr[34011]= -2015345591;
assign addr[34012]= -1987655498;
assign addr[34013]= -1957443913;
assign addr[34014]= -1924749160;
assign addr[34015]= -1889612716;
assign addr[34016]= -1852079154;
assign addr[34017]= -1812196087;
assign addr[34018]= -1770014111;
assign addr[34019]= -1725586737;
assign addr[34020]= -1678970324;
assign addr[34021]= -1630224009;
assign addr[34022]= -1579409630;
assign addr[34023]= -1526591649;
assign addr[34024]= -1471837070;
assign addr[34025]= -1415215352;
assign addr[34026]= -1356798326;
assign addr[34027]= -1296660098;
assign addr[34028]= -1234876957;
assign addr[34029]= -1171527280;
assign addr[34030]= -1106691431;
assign addr[34031]= -1040451659;
assign addr[34032]= -972891995;
assign addr[34033]= -904098143;
assign addr[34034]= -834157373;
assign addr[34035]= -763158411;
assign addr[34036]= -691191324;
assign addr[34037]= -618347408;
assign addr[34038]= -544719071;
assign addr[34039]= -470399716;
assign addr[34040]= -395483624;
assign addr[34041]= -320065829;
assign addr[34042]= -244242007;
assign addr[34043]= -168108346;
assign addr[34044]= -91761426;
assign addr[34045]= -15298099;
assign addr[34046]= 61184634;
assign addr[34047]= 137589750;
assign addr[34048]= 213820322;
assign addr[34049]= 289779648;
assign addr[34050]= 365371365;
assign addr[34051]= 440499581;
assign addr[34052]= 515068990;
assign addr[34053]= 588984994;
assign addr[34054]= 662153826;
assign addr[34055]= 734482665;
assign addr[34056]= 805879757;
assign addr[34057]= 876254528;
assign addr[34058]= 945517704;
assign addr[34059]= 1013581418;
assign addr[34060]= 1080359326;
assign addr[34061]= 1145766716;
assign addr[34062]= 1209720613;
assign addr[34063]= 1272139887;
assign addr[34064]= 1332945355;
assign addr[34065]= 1392059879;
assign addr[34066]= 1449408469;
assign addr[34067]= 1504918373;
assign addr[34068]= 1558519173;
assign addr[34069]= 1610142873;
assign addr[34070]= 1659723983;
assign addr[34071]= 1707199606;
assign addr[34072]= 1752509516;
assign addr[34073]= 1795596234;
assign addr[34074]= 1836405100;
assign addr[34075]= 1874884346;
assign addr[34076]= 1910985158;
assign addr[34077]= 1944661739;
assign addr[34078]= 1975871368;
assign addr[34079]= 2004574453;
assign addr[34080]= 2030734582;
assign addr[34081]= 2054318569;
assign addr[34082]= 2075296495;
assign addr[34083]= 2093641749;
assign addr[34084]= 2109331059;
assign addr[34085]= 2122344521;
assign addr[34086]= 2132665626;
assign addr[34087]= 2140281282;
assign addr[34088]= 2145181827;
assign addr[34089]= 2147361045;
assign addr[34090]= 2146816171;
assign addr[34091]= 2143547897;
assign addr[34092]= 2137560369;
assign addr[34093]= 2128861181;
assign addr[34094]= 2117461370;
assign addr[34095]= 2103375398;
assign addr[34096]= 2086621133;
assign addr[34097]= 2067219829;
assign addr[34098]= 2045196100;
assign addr[34099]= 2020577882;
assign addr[34100]= 1993396407;
assign addr[34101]= 1963686155;
assign addr[34102]= 1931484818;
assign addr[34103]= 1896833245;
assign addr[34104]= 1859775393;
assign addr[34105]= 1820358275;
assign addr[34106]= 1778631892;
assign addr[34107]= 1734649179;
assign addr[34108]= 1688465931;
assign addr[34109]= 1640140734;
assign addr[34110]= 1589734894;
assign addr[34111]= 1537312353;
assign addr[34112]= 1482939614;
assign addr[34113]= 1426685652;
assign addr[34114]= 1368621831;
assign addr[34115]= 1308821808;
assign addr[34116]= 1247361445;
assign addr[34117]= 1184318708;
assign addr[34118]= 1119773573;
assign addr[34119]= 1053807919;
assign addr[34120]= 986505429;
assign addr[34121]= 917951481;
assign addr[34122]= 848233042;
assign addr[34123]= 777438554;
assign addr[34124]= 705657826;
assign addr[34125]= 632981917;
assign addr[34126]= 559503022;
assign addr[34127]= 485314355;
assign addr[34128]= 410510029;
assign addr[34129]= 335184940;
assign addr[34130]= 259434643;
assign addr[34131]= 183355234;
assign addr[34132]= 107043224;
assign addr[34133]= 30595422;
assign addr[34134]= -45891193;
assign addr[34135]= -122319591;
assign addr[34136]= -198592817;
assign addr[34137]= -274614114;
assign addr[34138]= -350287041;
assign addr[34139]= -425515602;
assign addr[34140]= -500204365;
assign addr[34141]= -574258580;
assign addr[34142]= -647584304;
assign addr[34143]= -720088517;
assign addr[34144]= -791679244;
assign addr[34145]= -862265664;
assign addr[34146]= -931758235;
assign addr[34147]= -1000068799;
assign addr[34148]= -1067110699;
assign addr[34149]= -1132798888;
assign addr[34150]= -1197050035;
assign addr[34151]= -1259782632;
assign addr[34152]= -1320917099;
assign addr[34153]= -1380375881;
assign addr[34154]= -1438083551;
assign addr[34155]= -1493966902;
assign addr[34156]= -1547955041;
assign addr[34157]= -1599979481;
assign addr[34158]= -1649974225;
assign addr[34159]= -1697875851;
assign addr[34160]= -1743623590;
assign addr[34161]= -1787159411;
assign addr[34162]= -1828428082;
assign addr[34163]= -1867377253;
assign addr[34164]= -1903957513;
assign addr[34165]= -1938122457;
assign addr[34166]= -1969828744;
assign addr[34167]= -1999036154;
assign addr[34168]= -2025707632;
assign addr[34169]= -2049809346;
assign addr[34170]= -2071310720;
assign addr[34171]= -2090184478;
assign addr[34172]= -2106406677;
assign addr[34173]= -2119956737;
assign addr[34174]= -2130817471;
assign addr[34175]= -2138975100;
assign addr[34176]= -2144419275;
assign addr[34177]= -2147143090;
assign addr[34178]= -2147143090;
assign addr[34179]= -2144419275;
assign addr[34180]= -2138975100;
assign addr[34181]= -2130817471;
assign addr[34182]= -2119956737;
assign addr[34183]= -2106406677;
assign addr[34184]= -2090184478;
assign addr[34185]= -2071310720;
assign addr[34186]= -2049809346;
assign addr[34187]= -2025707632;
assign addr[34188]= -1999036154;
assign addr[34189]= -1969828744;
assign addr[34190]= -1938122457;
assign addr[34191]= -1903957513;
assign addr[34192]= -1867377253;
assign addr[34193]= -1828428082;
assign addr[34194]= -1787159411;
assign addr[34195]= -1743623590;
assign addr[34196]= -1697875851;
assign addr[34197]= -1649974225;
assign addr[34198]= -1599979481;
assign addr[34199]= -1547955041;
assign addr[34200]= -1493966902;
assign addr[34201]= -1438083551;
assign addr[34202]= -1380375881;
assign addr[34203]= -1320917099;
assign addr[34204]= -1259782632;
assign addr[34205]= -1197050035;
assign addr[34206]= -1132798888;
assign addr[34207]= -1067110699;
assign addr[34208]= -1000068799;
assign addr[34209]= -931758235;
assign addr[34210]= -862265664;
assign addr[34211]= -791679244;
assign addr[34212]= -720088517;
assign addr[34213]= -647584304;
assign addr[34214]= -574258580;
assign addr[34215]= -500204365;
assign addr[34216]= -425515602;
assign addr[34217]= -350287041;
assign addr[34218]= -274614114;
assign addr[34219]= -198592817;
assign addr[34220]= -122319591;
assign addr[34221]= -45891193;
assign addr[34222]= 30595422;
assign addr[34223]= 107043224;
assign addr[34224]= 183355234;
assign addr[34225]= 259434643;
assign addr[34226]= 335184940;
assign addr[34227]= 410510029;
assign addr[34228]= 485314355;
assign addr[34229]= 559503022;
assign addr[34230]= 632981917;
assign addr[34231]= 705657826;
assign addr[34232]= 777438554;
assign addr[34233]= 848233042;
assign addr[34234]= 917951481;
assign addr[34235]= 986505429;
assign addr[34236]= 1053807919;
assign addr[34237]= 1119773573;
assign addr[34238]= 1184318708;
assign addr[34239]= 1247361445;
assign addr[34240]= 1308821808;
assign addr[34241]= 1368621831;
assign addr[34242]= 1426685652;
assign addr[34243]= 1482939614;
assign addr[34244]= 1537312353;
assign addr[34245]= 1589734894;
assign addr[34246]= 1640140734;
assign addr[34247]= 1688465931;
assign addr[34248]= 1734649179;
assign addr[34249]= 1778631892;
assign addr[34250]= 1820358275;
assign addr[34251]= 1859775393;
assign addr[34252]= 1896833245;
assign addr[34253]= 1931484818;
assign addr[34254]= 1963686155;
assign addr[34255]= 1993396407;
assign addr[34256]= 2020577882;
assign addr[34257]= 2045196100;
assign addr[34258]= 2067219829;
assign addr[34259]= 2086621133;
assign addr[34260]= 2103375398;
assign addr[34261]= 2117461370;
assign addr[34262]= 2128861181;
assign addr[34263]= 2137560369;
assign addr[34264]= 2143547897;
assign addr[34265]= 2146816171;
assign addr[34266]= 2147361045;
assign addr[34267]= 2145181827;
assign addr[34268]= 2140281282;
assign addr[34269]= 2132665626;
assign addr[34270]= 2122344521;
assign addr[34271]= 2109331059;
assign addr[34272]= 2093641749;
assign addr[34273]= 2075296495;
assign addr[34274]= 2054318569;
assign addr[34275]= 2030734582;
assign addr[34276]= 2004574453;
assign addr[34277]= 1975871368;
assign addr[34278]= 1944661739;
assign addr[34279]= 1910985158;
assign addr[34280]= 1874884346;
assign addr[34281]= 1836405100;
assign addr[34282]= 1795596234;
assign addr[34283]= 1752509516;
assign addr[34284]= 1707199606;
assign addr[34285]= 1659723983;
assign addr[34286]= 1610142873;
assign addr[34287]= 1558519173;
assign addr[34288]= 1504918373;
assign addr[34289]= 1449408469;
assign addr[34290]= 1392059879;
assign addr[34291]= 1332945355;
assign addr[34292]= 1272139887;
assign addr[34293]= 1209720613;
assign addr[34294]= 1145766716;
assign addr[34295]= 1080359326;
assign addr[34296]= 1013581418;
assign addr[34297]= 945517704;
assign addr[34298]= 876254528;
assign addr[34299]= 805879757;
assign addr[34300]= 734482665;
assign addr[34301]= 662153826;
assign addr[34302]= 588984994;
assign addr[34303]= 515068990;
assign addr[34304]= 440499581;
assign addr[34305]= 365371365;
assign addr[34306]= 289779648;
assign addr[34307]= 213820322;
assign addr[34308]= 137589750;
assign addr[34309]= 61184634;
assign addr[34310]= -15298099;
assign addr[34311]= -91761426;
assign addr[34312]= -168108346;
assign addr[34313]= -244242007;
assign addr[34314]= -320065829;
assign addr[34315]= -395483624;
assign addr[34316]= -470399716;
assign addr[34317]= -544719071;
assign addr[34318]= -618347408;
assign addr[34319]= -691191324;
assign addr[34320]= -763158411;
assign addr[34321]= -834157373;
assign addr[34322]= -904098143;
assign addr[34323]= -972891995;
assign addr[34324]= -1040451659;
assign addr[34325]= -1106691431;
assign addr[34326]= -1171527280;
assign addr[34327]= -1234876957;
assign addr[34328]= -1296660098;
assign addr[34329]= -1356798326;
assign addr[34330]= -1415215352;
assign addr[34331]= -1471837070;
assign addr[34332]= -1526591649;
assign addr[34333]= -1579409630;
assign addr[34334]= -1630224009;
assign addr[34335]= -1678970324;
assign addr[34336]= -1725586737;
assign addr[34337]= -1770014111;
assign addr[34338]= -1812196087;
assign addr[34339]= -1852079154;
assign addr[34340]= -1889612716;
assign addr[34341]= -1924749160;
assign addr[34342]= -1957443913;
assign addr[34343]= -1987655498;
assign addr[34344]= -2015345591;
assign addr[34345]= -2040479063;
assign addr[34346]= -2063024031;
assign addr[34347]= -2082951896;
assign addr[34348]= -2100237377;
assign addr[34349]= -2114858546;
assign addr[34350]= -2126796855;
assign addr[34351]= -2136037160;
assign addr[34352]= -2142567738;
assign addr[34353]= -2146380306;
assign addr[34354]= -2147470025;
assign addr[34355]= -2145835515;
assign addr[34356]= -2141478848;
assign addr[34357]= -2134405552;
assign addr[34358]= -2124624598;
assign addr[34359]= -2112148396;
assign addr[34360]= -2096992772;
assign addr[34361]= -2079176953;
assign addr[34362]= -2058723538;
assign addr[34363]= -2035658475;
assign addr[34364]= -2010011024;
assign addr[34365]= -1981813720;
assign addr[34366]= -1951102334;
assign addr[34367]= -1917915825;
assign addr[34368]= -1882296293;
assign addr[34369]= -1844288924;
assign addr[34370]= -1803941934;
assign addr[34371]= -1761306505;
assign addr[34372]= -1716436725;
assign addr[34373]= -1669389513;
assign addr[34374]= -1620224553;
assign addr[34375]= -1569004214;
assign addr[34376]= -1515793473;
assign addr[34377]= -1460659832;
assign addr[34378]= -1403673233;
assign addr[34379]= -1344905966;
assign addr[34380]= -1284432584;
assign addr[34381]= -1222329801;
assign addr[34382]= -1158676398;
assign addr[34383]= -1093553126;
assign addr[34384]= -1027042599;
assign addr[34385]= -959229189;
assign addr[34386]= -890198924;
assign addr[34387]= -820039373;
assign addr[34388]= -748839539;
assign addr[34389]= -676689746;
assign addr[34390]= -603681519;
assign addr[34391]= -529907477;
assign addr[34392]= -455461206;
assign addr[34393]= -380437148;
assign addr[34394]= -304930476;
assign addr[34395]= -229036977;
assign addr[34396]= -152852926;
assign addr[34397]= -76474970;
assign addr[34398]= 0;
assign addr[34399]= 76474970;
assign addr[34400]= 152852926;
assign addr[34401]= 229036977;
assign addr[34402]= 304930476;
assign addr[34403]= 380437148;
assign addr[34404]= 455461206;
assign addr[34405]= 529907477;
assign addr[34406]= 603681519;
assign addr[34407]= 676689746;
assign addr[34408]= 748839539;
assign addr[34409]= 820039373;
assign addr[34410]= 890198924;
assign addr[34411]= 959229189;
assign addr[34412]= 1027042599;
assign addr[34413]= 1093553126;
assign addr[34414]= 1158676398;
assign addr[34415]= 1222329801;
assign addr[34416]= 1284432584;
assign addr[34417]= 1344905966;
assign addr[34418]= 1403673233;
assign addr[34419]= 1460659832;
assign addr[34420]= 1515793473;
assign addr[34421]= 1569004214;
assign addr[34422]= 1620224553;
assign addr[34423]= 1669389513;
assign addr[34424]= 1716436725;
assign addr[34425]= 1761306505;
assign addr[34426]= 1803941934;
assign addr[34427]= 1844288924;
assign addr[34428]= 1882296293;
assign addr[34429]= 1917915825;
assign addr[34430]= 1951102334;
assign addr[34431]= 1981813720;
assign addr[34432]= 2010011024;
assign addr[34433]= 2035658475;
assign addr[34434]= 2058723538;
assign addr[34435]= 2079176953;
assign addr[34436]= 2096992772;
assign addr[34437]= 2112148396;
assign addr[34438]= 2124624598;
assign addr[34439]= 2134405552;
assign addr[34440]= 2141478848;
assign addr[34441]= 2145835515;
assign addr[34442]= 2147470025;
assign addr[34443]= 2146380306;
assign addr[34444]= 2142567738;
assign addr[34445]= 2136037160;
assign addr[34446]= 2126796855;
assign addr[34447]= 2114858546;
assign addr[34448]= 2100237377;
assign addr[34449]= 2082951896;
assign addr[34450]= 2063024031;
assign addr[34451]= 2040479063;
assign addr[34452]= 2015345591;
assign addr[34453]= 1987655498;
assign addr[34454]= 1957443913;
assign addr[34455]= 1924749160;
assign addr[34456]= 1889612716;
assign addr[34457]= 1852079154;
assign addr[34458]= 1812196087;
assign addr[34459]= 1770014111;
assign addr[34460]= 1725586737;
assign addr[34461]= 1678970324;
assign addr[34462]= 1630224009;
assign addr[34463]= 1579409630;
assign addr[34464]= 1526591649;
assign addr[34465]= 1471837070;
assign addr[34466]= 1415215352;
assign addr[34467]= 1356798326;
assign addr[34468]= 1296660098;
assign addr[34469]= 1234876957;
assign addr[34470]= 1171527280;
assign addr[34471]= 1106691431;
assign addr[34472]= 1040451659;
assign addr[34473]= 972891995;
assign addr[34474]= 904098143;
assign addr[34475]= 834157373;
assign addr[34476]= 763158411;
assign addr[34477]= 691191324;
assign addr[34478]= 618347408;
assign addr[34479]= 544719071;
assign addr[34480]= 470399716;
assign addr[34481]= 395483624;
assign addr[34482]= 320065829;
assign addr[34483]= 244242007;
assign addr[34484]= 168108346;
assign addr[34485]= 91761426;
assign addr[34486]= 15298099;
assign addr[34487]= -61184634;
assign addr[34488]= -137589750;
assign addr[34489]= -213820322;
assign addr[34490]= -289779648;
assign addr[34491]= -365371365;
assign addr[34492]= -440499581;
assign addr[34493]= -515068990;
assign addr[34494]= -588984994;
assign addr[34495]= -662153826;
assign addr[34496]= -734482665;
assign addr[34497]= -805879757;
assign addr[34498]= -876254528;
assign addr[34499]= -945517704;
assign addr[34500]= -1013581418;
assign addr[34501]= -1080359326;
assign addr[34502]= -1145766716;
assign addr[34503]= -1209720613;
assign addr[34504]= -1272139887;
assign addr[34505]= -1332945355;
assign addr[34506]= -1392059879;
assign addr[34507]= -1449408469;
assign addr[34508]= -1504918373;
assign addr[34509]= -1558519173;
assign addr[34510]= -1610142873;
assign addr[34511]= -1659723983;
assign addr[34512]= -1707199606;
assign addr[34513]= -1752509516;
assign addr[34514]= -1795596234;
assign addr[34515]= -1836405100;
assign addr[34516]= -1874884346;
assign addr[34517]= -1910985158;
assign addr[34518]= -1944661739;
assign addr[34519]= -1975871368;
assign addr[34520]= -2004574453;
assign addr[34521]= -2030734582;
assign addr[34522]= -2054318569;
assign addr[34523]= -2075296495;
assign addr[34524]= -2093641749;
assign addr[34525]= -2109331059;
assign addr[34526]= -2122344521;
assign addr[34527]= -2132665626;
assign addr[34528]= -2140281282;
assign addr[34529]= -2145181827;
assign addr[34530]= -2147361045;
assign addr[34531]= -2146816171;
assign addr[34532]= -2143547897;
assign addr[34533]= -2137560369;
assign addr[34534]= -2128861181;
assign addr[34535]= -2117461370;
assign addr[34536]= -2103375398;
assign addr[34537]= -2086621133;
assign addr[34538]= -2067219829;
assign addr[34539]= -2045196100;
assign addr[34540]= -2020577882;
assign addr[34541]= -1993396407;
assign addr[34542]= -1963686155;
assign addr[34543]= -1931484818;
assign addr[34544]= -1896833245;
assign addr[34545]= -1859775393;
assign addr[34546]= -1820358275;
assign addr[34547]= -1778631892;
assign addr[34548]= -1734649179;
assign addr[34549]= -1688465931;
assign addr[34550]= -1640140734;
assign addr[34551]= -1589734894;
assign addr[34552]= -1537312353;
assign addr[34553]= -1482939614;
assign addr[34554]= -1426685652;
assign addr[34555]= -1368621831;
assign addr[34556]= -1308821808;
assign addr[34557]= -1247361445;
assign addr[34558]= -1184318708;
assign addr[34559]= -1119773573;
assign addr[34560]= -1053807919;
assign addr[34561]= -986505429;
assign addr[34562]= -917951481;
assign addr[34563]= -848233042;
assign addr[34564]= -777438554;
assign addr[34565]= -705657826;
assign addr[34566]= -632981917;
assign addr[34567]= -559503022;
assign addr[34568]= -485314355;
assign addr[34569]= -410510029;
assign addr[34570]= -335184940;
assign addr[34571]= -259434643;
assign addr[34572]= -183355234;
assign addr[34573]= -107043224;
assign addr[34574]= -30595422;
assign addr[34575]= 45891193;
assign addr[34576]= 122319591;
assign addr[34577]= 198592817;
assign addr[34578]= 274614114;
assign addr[34579]= 350287041;
assign addr[34580]= 425515602;
assign addr[34581]= 500204365;
assign addr[34582]= 574258580;
assign addr[34583]= 647584304;
assign addr[34584]= 720088517;
assign addr[34585]= 791679244;
assign addr[34586]= 862265664;
assign addr[34587]= 931758235;
assign addr[34588]= 1000068799;
assign addr[34589]= 1067110699;
assign addr[34590]= 1132798888;
assign addr[34591]= 1197050035;
assign addr[34592]= 1259782632;
assign addr[34593]= 1320917099;
assign addr[34594]= 1380375881;
assign addr[34595]= 1438083551;
assign addr[34596]= 1493966902;
assign addr[34597]= 1547955041;
assign addr[34598]= 1599979481;
assign addr[34599]= 1649974225;
assign addr[34600]= 1697875851;
assign addr[34601]= 1743623590;
assign addr[34602]= 1787159411;
assign addr[34603]= 1828428082;
assign addr[34604]= 1867377253;
assign addr[34605]= 1903957513;
assign addr[34606]= 1938122457;
assign addr[34607]= 1969828744;
assign addr[34608]= 1999036154;
assign addr[34609]= 2025707632;
assign addr[34610]= 2049809346;
assign addr[34611]= 2071310720;
assign addr[34612]= 2090184478;
assign addr[34613]= 2106406677;
assign addr[34614]= 2119956737;
assign addr[34615]= 2130817471;
assign addr[34616]= 2138975100;
assign addr[34617]= 2144419275;
assign addr[34618]= 2147143090;
assign addr[34619]= 2147143090;
assign addr[34620]= 2144419275;
assign addr[34621]= 2138975100;
assign addr[34622]= 2130817471;
assign addr[34623]= 2119956737;
assign addr[34624]= 2106406677;
assign addr[34625]= 2090184478;
assign addr[34626]= 2071310720;
assign addr[34627]= 2049809346;
assign addr[34628]= 2025707632;
assign addr[34629]= 1999036154;
assign addr[34630]= 1969828744;
assign addr[34631]= 1938122457;
assign addr[34632]= 1903957513;
assign addr[34633]= 1867377253;
assign addr[34634]= 1828428082;
assign addr[34635]= 1787159411;
assign addr[34636]= 1743623590;
assign addr[34637]= 1697875851;
assign addr[34638]= 1649974225;
assign addr[34639]= 1599979481;
assign addr[34640]= 1547955041;
assign addr[34641]= 1493966902;
assign addr[34642]= 1438083551;
assign addr[34643]= 1380375881;
assign addr[34644]= 1320917099;
assign addr[34645]= 1259782632;
assign addr[34646]= 1197050035;
assign addr[34647]= 1132798888;
assign addr[34648]= 1067110699;
assign addr[34649]= 1000068799;
assign addr[34650]= 931758235;
assign addr[34651]= 862265664;
assign addr[34652]= 791679244;
assign addr[34653]= 720088517;
assign addr[34654]= 647584304;
assign addr[34655]= 574258580;
assign addr[34656]= 500204365;
assign addr[34657]= 425515602;
assign addr[34658]= 350287041;
assign addr[34659]= 274614114;
assign addr[34660]= 198592817;
assign addr[34661]= 122319591;
assign addr[34662]= 45891193;
assign addr[34663]= -30595422;
assign addr[34664]= -107043224;
assign addr[34665]= -183355234;
assign addr[34666]= -259434643;
assign addr[34667]= -335184940;
assign addr[34668]= -410510029;
assign addr[34669]= -485314355;
assign addr[34670]= -559503022;
assign addr[34671]= -632981917;
assign addr[34672]= -705657826;
assign addr[34673]= -777438554;
assign addr[34674]= -848233042;
assign addr[34675]= -917951481;
assign addr[34676]= -986505429;
assign addr[34677]= -1053807919;
assign addr[34678]= -1119773573;
assign addr[34679]= -1184318708;
assign addr[34680]= -1247361445;
assign addr[34681]= -1308821808;
assign addr[34682]= -1368621831;
assign addr[34683]= -1426685652;
assign addr[34684]= -1482939614;
assign addr[34685]= -1537312353;
assign addr[34686]= -1589734894;
assign addr[34687]= -1640140734;
assign addr[34688]= -1688465931;
assign addr[34689]= -1734649179;
assign addr[34690]= -1778631892;
assign addr[34691]= -1820358275;
assign addr[34692]= -1859775393;
assign addr[34693]= -1896833245;
assign addr[34694]= -1931484818;
assign addr[34695]= -1963686155;
assign addr[34696]= -1993396407;
assign addr[34697]= -2020577882;
assign addr[34698]= -2045196100;
assign addr[34699]= -2067219829;
assign addr[34700]= -2086621133;
assign addr[34701]= -2103375398;
assign addr[34702]= -2117461370;
assign addr[34703]= -2128861181;
assign addr[34704]= -2137560369;
assign addr[34705]= -2143547897;
assign addr[34706]= -2146816171;
assign addr[34707]= -2147361045;
assign addr[34708]= -2145181827;
assign addr[34709]= -2140281282;
assign addr[34710]= -2132665626;
assign addr[34711]= -2122344521;
assign addr[34712]= -2109331059;
assign addr[34713]= -2093641749;
assign addr[34714]= -2075296495;
assign addr[34715]= -2054318569;
assign addr[34716]= -2030734582;
assign addr[34717]= -2004574453;
assign addr[34718]= -1975871368;
assign addr[34719]= -1944661739;
assign addr[34720]= -1910985158;
assign addr[34721]= -1874884346;
assign addr[34722]= -1836405100;
assign addr[34723]= -1795596234;
assign addr[34724]= -1752509516;
assign addr[34725]= -1707199606;
assign addr[34726]= -1659723983;
assign addr[34727]= -1610142873;
assign addr[34728]= -1558519173;
assign addr[34729]= -1504918373;
assign addr[34730]= -1449408469;
assign addr[34731]= -1392059879;
assign addr[34732]= -1332945355;
assign addr[34733]= -1272139887;
assign addr[34734]= -1209720613;
assign addr[34735]= -1145766716;
assign addr[34736]= -1080359326;
assign addr[34737]= -1013581418;
assign addr[34738]= -945517704;
assign addr[34739]= -876254528;
assign addr[34740]= -805879757;
assign addr[34741]= -734482665;
assign addr[34742]= -662153826;
assign addr[34743]= -588984994;
assign addr[34744]= -515068990;
assign addr[34745]= -440499581;
assign addr[34746]= -365371365;
assign addr[34747]= -289779648;
assign addr[34748]= -213820322;
assign addr[34749]= -137589750;
assign addr[34750]= -61184634;
assign addr[34751]= 15298099;
assign addr[34752]= 91761426;
assign addr[34753]= 168108346;
assign addr[34754]= 244242007;
assign addr[34755]= 320065829;
assign addr[34756]= 395483624;
assign addr[34757]= 470399716;
assign addr[34758]= 544719071;
assign addr[34759]= 618347408;
assign addr[34760]= 691191324;
assign addr[34761]= 763158411;
assign addr[34762]= 834157373;
assign addr[34763]= 904098143;
assign addr[34764]= 972891995;
assign addr[34765]= 1040451659;
assign addr[34766]= 1106691431;
assign addr[34767]= 1171527280;
assign addr[34768]= 1234876957;
assign addr[34769]= 1296660098;
assign addr[34770]= 1356798326;
assign addr[34771]= 1415215352;
assign addr[34772]= 1471837070;
assign addr[34773]= 1526591649;
assign addr[34774]= 1579409630;
assign addr[34775]= 1630224009;
assign addr[34776]= 1678970324;
assign addr[34777]= 1725586737;
assign addr[34778]= 1770014111;
assign addr[34779]= 1812196087;
assign addr[34780]= 1852079154;
assign addr[34781]= 1889612716;
assign addr[34782]= 1924749160;
assign addr[34783]= 1957443913;
assign addr[34784]= 1987655498;
assign addr[34785]= 2015345591;
assign addr[34786]= 2040479063;
assign addr[34787]= 2063024031;
assign addr[34788]= 2082951896;
assign addr[34789]= 2100237377;
assign addr[34790]= 2114858546;
assign addr[34791]= 2126796855;
assign addr[34792]= 2136037160;
assign addr[34793]= 2142567738;
assign addr[34794]= 2146380306;
assign addr[34795]= 2147470025;
assign addr[34796]= 2145835515;
assign addr[34797]= 2141478848;
assign addr[34798]= 2134405552;
assign addr[34799]= 2124624598;
assign addr[34800]= 2112148396;
assign addr[34801]= 2096992772;
assign addr[34802]= 2079176953;
assign addr[34803]= 2058723538;
assign addr[34804]= 2035658475;
assign addr[34805]= 2010011024;
assign addr[34806]= 1981813720;
assign addr[34807]= 1951102334;
assign addr[34808]= 1917915825;
assign addr[34809]= 1882296293;
assign addr[34810]= 1844288924;
assign addr[34811]= 1803941934;
assign addr[34812]= 1761306505;
assign addr[34813]= 1716436725;
assign addr[34814]= 1669389513;
assign addr[34815]= 1620224553;
assign addr[34816]= 1569004214;
assign addr[34817]= 1515793473;
assign addr[34818]= 1460659832;
assign addr[34819]= 1403673233;
assign addr[34820]= 1344905966;
assign addr[34821]= 1284432584;
assign addr[34822]= 1222329801;
assign addr[34823]= 1158676398;
assign addr[34824]= 1093553126;
assign addr[34825]= 1027042599;
assign addr[34826]= 959229189;
assign addr[34827]= 890198924;
assign addr[34828]= 820039373;
assign addr[34829]= 748839539;
assign addr[34830]= 676689746;
assign addr[34831]= 603681519;
assign addr[34832]= 529907477;
assign addr[34833]= 455461206;
assign addr[34834]= 380437148;
assign addr[34835]= 304930476;
assign addr[34836]= 229036977;
assign addr[34837]= 152852926;
assign addr[34838]= 76474970;
assign addr[34839]= 0;
assign addr[34840]= -76474970;
assign addr[34841]= -152852926;
assign addr[34842]= -229036977;
assign addr[34843]= -304930476;
assign addr[34844]= -380437148;
assign addr[34845]= -455461206;
assign addr[34846]= -529907477;
assign addr[34847]= -603681519;
assign addr[34848]= -676689746;
assign addr[34849]= -748839539;
assign addr[34850]= -820039373;
assign addr[34851]= -890198924;
assign addr[34852]= -959229189;
assign addr[34853]= -1027042599;
assign addr[34854]= -1093553126;
assign addr[34855]= -1158676398;
assign addr[34856]= -1222329801;
assign addr[34857]= -1284432584;
assign addr[34858]= -1344905966;
assign addr[34859]= -1403673233;
assign addr[34860]= -1460659832;
assign addr[34861]= -1515793473;
assign addr[34862]= -1569004214;
assign addr[34863]= -1620224553;
assign addr[34864]= -1669389513;
assign addr[34865]= -1716436725;
assign addr[34866]= -1761306505;
assign addr[34867]= -1803941934;
assign addr[34868]= -1844288924;
assign addr[34869]= -1882296293;
assign addr[34870]= -1917915825;
assign addr[34871]= -1951102334;
assign addr[34872]= -1981813720;
assign addr[34873]= -2010011024;
assign addr[34874]= -2035658475;
assign addr[34875]= -2058723538;
assign addr[34876]= -2079176953;
assign addr[34877]= -2096992772;
assign addr[34878]= -2112148396;
assign addr[34879]= -2124624598;
assign addr[34880]= -2134405552;
assign addr[34881]= -2141478848;
assign addr[34882]= -2145835515;
assign addr[34883]= -2147470025;
assign addr[34884]= -2146380306;
assign addr[34885]= -2142567738;
assign addr[34886]= -2136037160;
assign addr[34887]= -2126796855;
assign addr[34888]= -2114858546;
assign addr[34889]= -2100237377;
assign addr[34890]= -2082951896;
assign addr[34891]= -2063024031;
assign addr[34892]= -2040479063;
assign addr[34893]= -2015345591;
assign addr[34894]= -1987655498;
assign addr[34895]= -1957443913;
assign addr[34896]= -1924749160;
assign addr[34897]= -1889612716;
assign addr[34898]= -1852079154;
assign addr[34899]= -1812196087;
assign addr[34900]= -1770014111;
assign addr[34901]= -1725586737;
assign addr[34902]= -1678970324;
assign addr[34903]= -1630224009;
assign addr[34904]= -1579409630;
assign addr[34905]= -1526591649;
assign addr[34906]= -1471837070;
assign addr[34907]= -1415215352;
assign addr[34908]= -1356798326;
assign addr[34909]= -1296660098;
assign addr[34910]= -1234876957;
assign addr[34911]= -1171527280;
assign addr[34912]= -1106691431;
assign addr[34913]= -1040451659;
assign addr[34914]= -972891995;
assign addr[34915]= -904098143;
assign addr[34916]= -834157373;
assign addr[34917]= -763158411;
assign addr[34918]= -691191324;
assign addr[34919]= -618347408;
assign addr[34920]= -544719071;
assign addr[34921]= -470399716;
assign addr[34922]= -395483624;
assign addr[34923]= -320065829;
assign addr[34924]= -244242007;
assign addr[34925]= -168108346;
assign addr[34926]= -91761426;
assign addr[34927]= -15298099;
assign addr[34928]= 61184634;
assign addr[34929]= 137589750;
assign addr[34930]= 213820322;
assign addr[34931]= 289779648;
assign addr[34932]= 365371365;
assign addr[34933]= 440499581;
assign addr[34934]= 515068990;
assign addr[34935]= 588984994;
assign addr[34936]= 662153826;
assign addr[34937]= 734482665;
assign addr[34938]= 805879757;
assign addr[34939]= 876254528;
assign addr[34940]= 945517704;
assign addr[34941]= 1013581418;
assign addr[34942]= 1080359326;
assign addr[34943]= 1145766716;
assign addr[34944]= 1209720613;
assign addr[34945]= 1272139887;
assign addr[34946]= 1332945355;
assign addr[34947]= 1392059879;
assign addr[34948]= 1449408469;
assign addr[34949]= 1504918373;
assign addr[34950]= 1558519173;
assign addr[34951]= 1610142873;
assign addr[34952]= 1659723983;
assign addr[34953]= 1707199606;
assign addr[34954]= 1752509516;
assign addr[34955]= 1795596234;
assign addr[34956]= 1836405100;
assign addr[34957]= 1874884346;
assign addr[34958]= 1910985158;
assign addr[34959]= 1944661739;
assign addr[34960]= 1975871368;
assign addr[34961]= 2004574453;
assign addr[34962]= 2030734582;
assign addr[34963]= 2054318569;
assign addr[34964]= 2075296495;
assign addr[34965]= 2093641749;
assign addr[34966]= 2109331059;
assign addr[34967]= 2122344521;
assign addr[34968]= 2132665626;
assign addr[34969]= 2140281282;
assign addr[34970]= 2145181827;
assign addr[34971]= 2147361045;
assign addr[34972]= 2146816171;
assign addr[34973]= 2143547897;
assign addr[34974]= 2137560369;
assign addr[34975]= 2128861181;
assign addr[34976]= 2117461370;
assign addr[34977]= 2103375398;
assign addr[34978]= 2086621133;
assign addr[34979]= 2067219829;
assign addr[34980]= 2045196100;
assign addr[34981]= 2020577882;
assign addr[34982]= 1993396407;
assign addr[34983]= 1963686155;
assign addr[34984]= 1931484818;
assign addr[34985]= 1896833245;
assign addr[34986]= 1859775393;
assign addr[34987]= 1820358275;
assign addr[34988]= 1778631892;
assign addr[34989]= 1734649179;
assign addr[34990]= 1688465931;
assign addr[34991]= 1640140734;
assign addr[34992]= 1589734894;
assign addr[34993]= 1537312353;
assign addr[34994]= 1482939614;
assign addr[34995]= 1426685652;
assign addr[34996]= 1368621831;
assign addr[34997]= 1308821808;
assign addr[34998]= 1247361445;
assign addr[34999]= 1184318708;
assign addr[35000]= 1119773573;
assign addr[35001]= 1053807919;
assign addr[35002]= 986505429;
assign addr[35003]= 917951481;
assign addr[35004]= 848233042;
assign addr[35005]= 777438554;
assign addr[35006]= 705657826;
assign addr[35007]= 632981917;
assign addr[35008]= 559503022;
assign addr[35009]= 485314355;
assign addr[35010]= 410510029;
assign addr[35011]= 335184940;
assign addr[35012]= 259434643;
assign addr[35013]= 183355234;
assign addr[35014]= 107043224;
assign addr[35015]= 30595422;
assign addr[35016]= -45891193;
assign addr[35017]= -122319591;
assign addr[35018]= -198592817;
assign addr[35019]= -274614114;
assign addr[35020]= -350287041;
assign addr[35021]= -425515602;
assign addr[35022]= -500204365;
assign addr[35023]= -574258580;
assign addr[35024]= -647584304;
assign addr[35025]= -720088517;
assign addr[35026]= -791679244;
assign addr[35027]= -862265664;
assign addr[35028]= -931758235;
assign addr[35029]= -1000068799;
assign addr[35030]= -1067110699;
assign addr[35031]= -1132798888;
assign addr[35032]= -1197050035;
assign addr[35033]= -1259782632;
assign addr[35034]= -1320917099;
assign addr[35035]= -1380375881;
assign addr[35036]= -1438083551;
assign addr[35037]= -1493966902;
assign addr[35038]= -1547955041;
assign addr[35039]= -1599979481;
assign addr[35040]= -1649974225;
assign addr[35041]= -1697875851;
assign addr[35042]= -1743623590;
assign addr[35043]= -1787159411;
assign addr[35044]= -1828428082;
assign addr[35045]= -1867377253;
assign addr[35046]= -1903957513;
assign addr[35047]= -1938122457;
assign addr[35048]= -1969828744;
assign addr[35049]= -1999036154;
assign addr[35050]= -2025707632;
assign addr[35051]= -2049809346;
assign addr[35052]= -2071310720;
assign addr[35053]= -2090184478;
assign addr[35054]= -2106406677;
assign addr[35055]= -2119956737;
assign addr[35056]= -2130817471;
assign addr[35057]= -2138975100;
assign addr[35058]= -2144419275;
assign addr[35059]= -2147143090;
assign addr[35060]= -2147143090;
assign addr[35061]= -2144419275;
assign addr[35062]= -2138975100;
assign addr[35063]= -2130817471;
assign addr[35064]= -2119956737;
assign addr[35065]= -2106406677;
assign addr[35066]= -2090184478;
assign addr[35067]= -2071310720;
assign addr[35068]= -2049809346;
assign addr[35069]= -2025707632;
assign addr[35070]= -1999036154;
assign addr[35071]= -1969828744;
assign addr[35072]= -1938122457;
assign addr[35073]= -1903957513;
assign addr[35074]= -1867377253;
assign addr[35075]= -1828428082;
assign addr[35076]= -1787159411;
assign addr[35077]= -1743623590;
assign addr[35078]= -1697875851;
assign addr[35079]= -1649974225;
assign addr[35080]= -1599979481;
assign addr[35081]= -1547955041;
assign addr[35082]= -1493966902;
assign addr[35083]= -1438083551;
assign addr[35084]= -1380375881;
assign addr[35085]= -1320917099;
assign addr[35086]= -1259782632;
assign addr[35087]= -1197050035;
assign addr[35088]= -1132798888;
assign addr[35089]= -1067110699;
assign addr[35090]= -1000068799;
assign addr[35091]= -931758235;
assign addr[35092]= -862265664;
assign addr[35093]= -791679244;
assign addr[35094]= -720088517;
assign addr[35095]= -647584304;
assign addr[35096]= -574258580;
assign addr[35097]= -500204365;
assign addr[35098]= -425515602;
assign addr[35099]= -350287041;
assign addr[35100]= -274614114;
assign addr[35101]= -198592817;
assign addr[35102]= -122319591;
assign addr[35103]= -45891193;
assign addr[35104]= 30595422;
assign addr[35105]= 107043224;
assign addr[35106]= 183355234;
assign addr[35107]= 259434643;
assign addr[35108]= 335184940;
assign addr[35109]= 410510029;
assign addr[35110]= 485314355;
assign addr[35111]= 559503022;
assign addr[35112]= 632981917;
assign addr[35113]= 705657826;
assign addr[35114]= 777438554;
assign addr[35115]= 848233042;
assign addr[35116]= 917951481;
assign addr[35117]= 986505429;
assign addr[35118]= 1053807919;
assign addr[35119]= 1119773573;
assign addr[35120]= 1184318708;
assign addr[35121]= 1247361445;
assign addr[35122]= 1308821808;
assign addr[35123]= 1368621831;
assign addr[35124]= 1426685652;
assign addr[35125]= 1482939614;
assign addr[35126]= 1537312353;
assign addr[35127]= 1589734894;
assign addr[35128]= 1640140734;
assign addr[35129]= 1688465931;
assign addr[35130]= 1734649179;
assign addr[35131]= 1778631892;
assign addr[35132]= 1820358275;
assign addr[35133]= 1859775393;
assign addr[35134]= 1896833245;
assign addr[35135]= 1931484818;
assign addr[35136]= 1963686155;
assign addr[35137]= 1993396407;
assign addr[35138]= 2020577882;
assign addr[35139]= 2045196100;
assign addr[35140]= 2067219829;
assign addr[35141]= 2086621133;
assign addr[35142]= 2103375398;
assign addr[35143]= 2117461370;
assign addr[35144]= 2128861181;
assign addr[35145]= 2137560369;
assign addr[35146]= 2143547897;
assign addr[35147]= 2146816171;
assign addr[35148]= 2147361045;
assign addr[35149]= 2145181827;
assign addr[35150]= 2140281282;
assign addr[35151]= 2132665626;
assign addr[35152]= 2122344521;
assign addr[35153]= 2109331059;
assign addr[35154]= 2093641749;
assign addr[35155]= 2075296495;
assign addr[35156]= 2054318569;
assign addr[35157]= 2030734582;
assign addr[35158]= 2004574453;
assign addr[35159]= 1975871368;
assign addr[35160]= 1944661739;
assign addr[35161]= 1910985158;
assign addr[35162]= 1874884346;
assign addr[35163]= 1836405100;
assign addr[35164]= 1795596234;
assign addr[35165]= 1752509516;
assign addr[35166]= 1707199606;
assign addr[35167]= 1659723983;
assign addr[35168]= 1610142873;
assign addr[35169]= 1558519173;
assign addr[35170]= 1504918373;
assign addr[35171]= 1449408469;
assign addr[35172]= 1392059879;
assign addr[35173]= 1332945355;
assign addr[35174]= 1272139887;
assign addr[35175]= 1209720613;
assign addr[35176]= 1145766716;
assign addr[35177]= 1080359326;
assign addr[35178]= 1013581418;
assign addr[35179]= 945517704;
assign addr[35180]= 876254528;
assign addr[35181]= 805879757;
assign addr[35182]= 734482665;
assign addr[35183]= 662153826;
assign addr[35184]= 588984994;
assign addr[35185]= 515068990;
assign addr[35186]= 440499581;
assign addr[35187]= 365371365;
assign addr[35188]= 289779648;
assign addr[35189]= 213820322;
assign addr[35190]= 137589750;
assign addr[35191]= 61184634;
assign addr[35192]= -15298099;
assign addr[35193]= -91761426;
assign addr[35194]= -168108346;
assign addr[35195]= -244242007;
assign addr[35196]= -320065829;
assign addr[35197]= -395483624;
assign addr[35198]= -470399716;
assign addr[35199]= -544719071;
assign addr[35200]= -618347408;
assign addr[35201]= -691191324;
assign addr[35202]= -763158411;
assign addr[35203]= -834157373;
assign addr[35204]= -904098143;
assign addr[35205]= -972891995;
assign addr[35206]= -1040451659;
assign addr[35207]= -1106691431;
assign addr[35208]= -1171527280;
assign addr[35209]= -1234876957;
assign addr[35210]= -1296660098;
assign addr[35211]= -1356798326;
assign addr[35212]= -1415215352;
assign addr[35213]= -1471837070;
assign addr[35214]= -1526591649;
assign addr[35215]= -1579409630;
assign addr[35216]= -1630224009;
assign addr[35217]= -1678970324;
assign addr[35218]= -1725586737;
assign addr[35219]= -1770014111;
assign addr[35220]= -1812196087;
assign addr[35221]= -1852079154;
assign addr[35222]= -1889612716;
assign addr[35223]= -1924749160;
assign addr[35224]= -1957443913;
assign addr[35225]= -1987655498;
assign addr[35226]= -2015345591;
assign addr[35227]= -2040479063;
assign addr[35228]= -2063024031;
assign addr[35229]= -2082951896;
assign addr[35230]= -2100237377;
assign addr[35231]= -2114858546;
assign addr[35232]= -2126796855;
assign addr[35233]= -2136037160;
assign addr[35234]= -2142567738;
assign addr[35235]= -2146380306;
assign addr[35236]= -2147470025;
assign addr[35237]= -2145835515;
assign addr[35238]= -2141478848;
assign addr[35239]= -2134405552;
assign addr[35240]= -2124624598;
assign addr[35241]= -2112148396;
assign addr[35242]= -2096992772;
assign addr[35243]= -2079176953;
assign addr[35244]= -2058723538;
assign addr[35245]= -2035658475;
assign addr[35246]= -2010011024;
assign addr[35247]= -1981813720;
assign addr[35248]= -1951102334;
assign addr[35249]= -1917915825;
assign addr[35250]= -1882296293;
assign addr[35251]= -1844288924;
assign addr[35252]= -1803941934;
assign addr[35253]= -1761306505;
assign addr[35254]= -1716436725;
assign addr[35255]= -1669389513;
assign addr[35256]= -1620224553;
assign addr[35257]= -1569004214;
assign addr[35258]= -1515793473;
assign addr[35259]= -1460659832;
assign addr[35260]= -1403673233;
assign addr[35261]= -1344905966;
assign addr[35262]= -1284432584;
assign addr[35263]= -1222329801;
assign addr[35264]= -1158676398;
assign addr[35265]= -1093553126;
assign addr[35266]= -1027042599;
assign addr[35267]= -959229189;
assign addr[35268]= -890198924;
assign addr[35269]= -820039373;
assign addr[35270]= -748839539;
assign addr[35271]= -676689746;
assign addr[35272]= -603681519;
assign addr[35273]= -529907477;
assign addr[35274]= -455461206;
assign addr[35275]= -380437148;
assign addr[35276]= -304930476;
assign addr[35277]= -229036977;
assign addr[35278]= -152852926;
assign addr[35279]= -76474970;
assign addr[35280]= 0;
assign addr[35281]= 76474970;
assign addr[35282]= 152852926;
assign addr[35283]= 229036977;
assign addr[35284]= 304930476;
assign addr[35285]= 380437148;
assign addr[35286]= 455461206;
assign addr[35287]= 529907477;
assign addr[35288]= 603681519;
assign addr[35289]= 676689746;
assign addr[35290]= 748839539;
assign addr[35291]= 820039373;
assign addr[35292]= 890198924;
assign addr[35293]= 959229189;
assign addr[35294]= 1027042599;
assign addr[35295]= 1093553126;
assign addr[35296]= 1158676398;
assign addr[35297]= 1222329801;
assign addr[35298]= 1284432584;
assign addr[35299]= 1344905966;
assign addr[35300]= 1403673233;
assign addr[35301]= 1460659832;
assign addr[35302]= 1515793473;
assign addr[35303]= 1569004214;
assign addr[35304]= 1620224553;
assign addr[35305]= 1669389513;
assign addr[35306]= 1716436725;
assign addr[35307]= 1761306505;
assign addr[35308]= 1803941934;
assign addr[35309]= 1844288924;
assign addr[35310]= 1882296293;
assign addr[35311]= 1917915825;
assign addr[35312]= 1951102334;
assign addr[35313]= 1981813720;
assign addr[35314]= 2010011024;
assign addr[35315]= 2035658475;
assign addr[35316]= 2058723538;
assign addr[35317]= 2079176953;
assign addr[35318]= 2096992772;
assign addr[35319]= 2112148396;
assign addr[35320]= 2124624598;
assign addr[35321]= 2134405552;
assign addr[35322]= 2141478848;
assign addr[35323]= 2145835515;
assign addr[35324]= 2147470025;
assign addr[35325]= 2146380306;
assign addr[35326]= 2142567738;
assign addr[35327]= 2136037160;
assign addr[35328]= 2126796855;
assign addr[35329]= 2114858546;
assign addr[35330]= 2100237377;
assign addr[35331]= 2082951896;
assign addr[35332]= 2063024031;
assign addr[35333]= 2040479063;
assign addr[35334]= 2015345591;
assign addr[35335]= 1987655498;
assign addr[35336]= 1957443913;
assign addr[35337]= 1924749160;
assign addr[35338]= 1889612716;
assign addr[35339]= 1852079154;
assign addr[35340]= 1812196087;
assign addr[35341]= 1770014111;
assign addr[35342]= 1725586737;
assign addr[35343]= 1678970324;
assign addr[35344]= 1630224009;
assign addr[35345]= 1579409630;
assign addr[35346]= 1526591649;
assign addr[35347]= 1471837070;
assign addr[35348]= 1415215352;
assign addr[35349]= 1356798326;
assign addr[35350]= 1296660098;
assign addr[35351]= 1234876957;
assign addr[35352]= 1171527280;
assign addr[35353]= 1106691431;
assign addr[35354]= 1040451659;
assign addr[35355]= 972891995;
assign addr[35356]= 904098143;
assign addr[35357]= 834157373;
assign addr[35358]= 763158411;
assign addr[35359]= 691191324;
assign addr[35360]= 618347408;
assign addr[35361]= 544719071;
assign addr[35362]= 470399716;
assign addr[35363]= 395483624;
assign addr[35364]= 320065829;
assign addr[35365]= 244242007;
assign addr[35366]= 168108346;
assign addr[35367]= 91761426;
assign addr[35368]= 15298099;
assign addr[35369]= -61184634;
assign addr[35370]= -137589750;
assign addr[35371]= -213820322;
assign addr[35372]= -289779648;
assign addr[35373]= -365371365;
assign addr[35374]= -440499581;
assign addr[35375]= -515068990;
assign addr[35376]= -588984994;
assign addr[35377]= -662153826;
assign addr[35378]= -734482665;
assign addr[35379]= -805879757;
assign addr[35380]= -876254528;
assign addr[35381]= -945517704;
assign addr[35382]= -1013581418;
assign addr[35383]= -1080359326;
assign addr[35384]= -1145766716;
assign addr[35385]= -1209720613;
assign addr[35386]= -1272139887;
assign addr[35387]= -1332945355;
assign addr[35388]= -1392059879;
assign addr[35389]= -1449408469;
assign addr[35390]= -1504918373;
assign addr[35391]= -1558519173;
assign addr[35392]= -1610142873;
assign addr[35393]= -1659723983;
assign addr[35394]= -1707199606;
assign addr[35395]= -1752509516;
assign addr[35396]= -1795596234;
assign addr[35397]= -1836405100;
assign addr[35398]= -1874884346;
assign addr[35399]= -1910985158;
assign addr[35400]= -1944661739;
assign addr[35401]= -1975871368;
assign addr[35402]= -2004574453;
assign addr[35403]= -2030734582;
assign addr[35404]= -2054318569;
assign addr[35405]= -2075296495;
assign addr[35406]= -2093641749;
assign addr[35407]= -2109331059;
assign addr[35408]= -2122344521;
assign addr[35409]= -2132665626;
assign addr[35410]= -2140281282;
assign addr[35411]= -2145181827;
assign addr[35412]= -2147361045;
assign addr[35413]= -2146816171;
assign addr[35414]= -2143547897;
assign addr[35415]= -2137560369;
assign addr[35416]= -2128861181;
assign addr[35417]= -2117461370;
assign addr[35418]= -2103375398;
assign addr[35419]= -2086621133;
assign addr[35420]= -2067219829;
assign addr[35421]= -2045196100;
assign addr[35422]= -2020577882;
assign addr[35423]= -1993396407;
assign addr[35424]= -1963686155;
assign addr[35425]= -1931484818;
assign addr[35426]= -1896833245;
assign addr[35427]= -1859775393;
assign addr[35428]= -1820358275;
assign addr[35429]= -1778631892;
assign addr[35430]= -1734649179;
assign addr[35431]= -1688465931;
assign addr[35432]= -1640140734;
assign addr[35433]= -1589734894;
assign addr[35434]= -1537312353;
assign addr[35435]= -1482939614;
assign addr[35436]= -1426685652;
assign addr[35437]= -1368621831;
assign addr[35438]= -1308821808;
assign addr[35439]= -1247361445;
assign addr[35440]= -1184318708;
assign addr[35441]= -1119773573;
assign addr[35442]= -1053807919;
assign addr[35443]= -986505429;
assign addr[35444]= -917951481;
assign addr[35445]= -848233042;
assign addr[35446]= -777438554;
assign addr[35447]= -705657826;
assign addr[35448]= -632981917;
assign addr[35449]= -559503022;
assign addr[35450]= -485314355;
assign addr[35451]= -410510029;
assign addr[35452]= -335184940;
assign addr[35453]= -259434643;
assign addr[35454]= -183355234;
assign addr[35455]= -107043224;
assign addr[35456]= -30595422;
assign addr[35457]= 45891193;
assign addr[35458]= 122319591;
assign addr[35459]= 198592817;
assign addr[35460]= 274614114;
assign addr[35461]= 350287041;
assign addr[35462]= 425515602;
assign addr[35463]= 500204365;
assign addr[35464]= 574258580;
assign addr[35465]= 647584304;
assign addr[35466]= 720088517;
assign addr[35467]= 791679244;
assign addr[35468]= 862265664;
assign addr[35469]= 931758235;
assign addr[35470]= 1000068799;
assign addr[35471]= 1067110699;
assign addr[35472]= 1132798888;
assign addr[35473]= 1197050035;
assign addr[35474]= 1259782632;
assign addr[35475]= 1320917099;
assign addr[35476]= 1380375881;
assign addr[35477]= 1438083551;
assign addr[35478]= 1493966902;
assign addr[35479]= 1547955041;
assign addr[35480]= 1599979481;
assign addr[35481]= 1649974225;
assign addr[35482]= 1697875851;
assign addr[35483]= 1743623590;
assign addr[35484]= 1787159411;
assign addr[35485]= 1828428082;
assign addr[35486]= 1867377253;
assign addr[35487]= 1903957513;
assign addr[35488]= 1938122457;
assign addr[35489]= 1969828744;
assign addr[35490]= 1999036154;
assign addr[35491]= 2025707632;
assign addr[35492]= 2049809346;
assign addr[35493]= 2071310720;
assign addr[35494]= 2090184478;
assign addr[35495]= 2106406677;
assign addr[35496]= 2119956737;
assign addr[35497]= 2130817471;
assign addr[35498]= 2138975100;
assign addr[35499]= 2144419275;
assign addr[35500]= 2147143090;
assign addr[35501]= 2147143090;
assign addr[35502]= 2144419275;
assign addr[35503]= 2138975100;
assign addr[35504]= 2130817471;
assign addr[35505]= 2119956737;
assign addr[35506]= 2106406677;
assign addr[35507]= 2090184478;
assign addr[35508]= 2071310720;
assign addr[35509]= 2049809346;
assign addr[35510]= 2025707632;
assign addr[35511]= 1999036154;
assign addr[35512]= 1969828744;
assign addr[35513]= 1938122457;
assign addr[35514]= 1903957513;
assign addr[35515]= 1867377253;
assign addr[35516]= 1828428082;
assign addr[35517]= 1787159411;
assign addr[35518]= 1743623590;
assign addr[35519]= 1697875851;
assign addr[35520]= 1649974225;
assign addr[35521]= 1599979481;
assign addr[35522]= 1547955041;
assign addr[35523]= 1493966902;
assign addr[35524]= 1438083551;
assign addr[35525]= 1380375881;
assign addr[35526]= 1320917099;
assign addr[35527]= 1259782632;
assign addr[35528]= 1197050035;
assign addr[35529]= 1132798888;
assign addr[35530]= 1067110699;
assign addr[35531]= 1000068799;
assign addr[35532]= 931758235;
assign addr[35533]= 862265664;
assign addr[35534]= 791679244;
assign addr[35535]= 720088517;
assign addr[35536]= 647584304;
assign addr[35537]= 574258580;
assign addr[35538]= 500204365;
assign addr[35539]= 425515602;
assign addr[35540]= 350287041;
assign addr[35541]= 274614114;
assign addr[35542]= 198592817;
assign addr[35543]= 122319591;
assign addr[35544]= 45891193;
assign addr[35545]= -30595422;
assign addr[35546]= -107043224;
assign addr[35547]= -183355234;
assign addr[35548]= -259434643;
assign addr[35549]= -335184940;
assign addr[35550]= -410510029;
assign addr[35551]= -485314355;
assign addr[35552]= -559503022;
assign addr[35553]= -632981917;
assign addr[35554]= -705657826;
assign addr[35555]= -777438554;
assign addr[35556]= -848233042;
assign addr[35557]= -917951481;
assign addr[35558]= -986505429;
assign addr[35559]= -1053807919;
assign addr[35560]= -1119773573;
assign addr[35561]= -1184318708;
assign addr[35562]= -1247361445;
assign addr[35563]= -1308821808;
assign addr[35564]= -1368621831;
assign addr[35565]= -1426685652;
assign addr[35566]= -1482939614;
assign addr[35567]= -1537312353;
assign addr[35568]= -1589734894;
assign addr[35569]= -1640140734;
assign addr[35570]= -1688465931;
assign addr[35571]= -1734649179;
assign addr[35572]= -1778631892;
assign addr[35573]= -1820358275;
assign addr[35574]= -1859775393;
assign addr[35575]= -1896833245;
assign addr[35576]= -1931484818;
assign addr[35577]= -1963686155;
assign addr[35578]= -1993396407;
assign addr[35579]= -2020577882;
assign addr[35580]= -2045196100;
assign addr[35581]= -2067219829;
assign addr[35582]= -2086621133;
assign addr[35583]= -2103375398;
assign addr[35584]= -2117461370;
assign addr[35585]= -2128861181;
assign addr[35586]= -2137560369;
assign addr[35587]= -2143547897;
assign addr[35588]= -2146816171;
assign addr[35589]= -2147361045;
assign addr[35590]= -2145181827;
assign addr[35591]= -2140281282;
assign addr[35592]= -2132665626;
assign addr[35593]= -2122344521;
assign addr[35594]= -2109331059;
assign addr[35595]= -2093641749;
assign addr[35596]= -2075296495;
assign addr[35597]= -2054318569;
assign addr[35598]= -2030734582;
assign addr[35599]= -2004574453;
assign addr[35600]= -1975871368;
assign addr[35601]= -1944661739;
assign addr[35602]= -1910985158;
assign addr[35603]= -1874884346;
assign addr[35604]= -1836405100;
assign addr[35605]= -1795596234;
assign addr[35606]= -1752509516;
assign addr[35607]= -1707199606;
assign addr[35608]= -1659723983;
assign addr[35609]= -1610142873;
assign addr[35610]= -1558519173;
assign addr[35611]= -1504918373;
assign addr[35612]= -1449408469;
assign addr[35613]= -1392059879;
assign addr[35614]= -1332945355;
assign addr[35615]= -1272139887;
assign addr[35616]= -1209720613;
assign addr[35617]= -1145766716;
assign addr[35618]= -1080359326;
assign addr[35619]= -1013581418;
assign addr[35620]= -945517704;
assign addr[35621]= -876254528;
assign addr[35622]= -805879757;
assign addr[35623]= -734482665;
assign addr[35624]= -662153826;
assign addr[35625]= -588984994;
assign addr[35626]= -515068990;
assign addr[35627]= -440499581;
assign addr[35628]= -365371365;
assign addr[35629]= -289779648;
assign addr[35630]= -213820322;
assign addr[35631]= -137589750;
assign addr[35632]= -61184634;
assign addr[35633]= 15298099;
assign addr[35634]= 91761426;
assign addr[35635]= 168108346;
assign addr[35636]= 244242007;
assign addr[35637]= 320065829;
assign addr[35638]= 395483624;
assign addr[35639]= 470399716;
assign addr[35640]= 544719071;
assign addr[35641]= 618347408;
assign addr[35642]= 691191324;
assign addr[35643]= 763158411;
assign addr[35644]= 834157373;
assign addr[35645]= 904098143;
assign addr[35646]= 972891995;
assign addr[35647]= 1040451659;
assign addr[35648]= 1106691431;
assign addr[35649]= 1171527280;
assign addr[35650]= 1234876957;
assign addr[35651]= 1296660098;
assign addr[35652]= 1356798326;
assign addr[35653]= 1415215352;
assign addr[35654]= 1471837070;
assign addr[35655]= 1526591649;
assign addr[35656]= 1579409630;
assign addr[35657]= 1630224009;
assign addr[35658]= 1678970324;
assign addr[35659]= 1725586737;
assign addr[35660]= 1770014111;
assign addr[35661]= 1812196087;
assign addr[35662]= 1852079154;
assign addr[35663]= 1889612716;
assign addr[35664]= 1924749160;
assign addr[35665]= 1957443913;
assign addr[35666]= 1987655498;
assign addr[35667]= 2015345591;
assign addr[35668]= 2040479063;
assign addr[35669]= 2063024031;
assign addr[35670]= 2082951896;
assign addr[35671]= 2100237377;
assign addr[35672]= 2114858546;
assign addr[35673]= 2126796855;
assign addr[35674]= 2136037160;
assign addr[35675]= 2142567738;
assign addr[35676]= 2146380306;
assign addr[35677]= 2147470025;
assign addr[35678]= 2145835515;
assign addr[35679]= 2141478848;
assign addr[35680]= 2134405552;
assign addr[35681]= 2124624598;
assign addr[35682]= 2112148396;
assign addr[35683]= 2096992772;
assign addr[35684]= 2079176953;
assign addr[35685]= 2058723538;
assign addr[35686]= 2035658475;
assign addr[35687]= 2010011024;
assign addr[35688]= 1981813720;
assign addr[35689]= 1951102334;
assign addr[35690]= 1917915825;
assign addr[35691]= 1882296293;
assign addr[35692]= 1844288924;
assign addr[35693]= 1803941934;
assign addr[35694]= 1761306505;
assign addr[35695]= 1716436725;
assign addr[35696]= 1669389513;
assign addr[35697]= 1620224553;
assign addr[35698]= 1569004214;
assign addr[35699]= 1515793473;
assign addr[35700]= 1460659832;
assign addr[35701]= 1403673233;
assign addr[35702]= 1344905966;
assign addr[35703]= 1284432584;
assign addr[35704]= 1222329801;
assign addr[35705]= 1158676398;
assign addr[35706]= 1093553126;
assign addr[35707]= 1027042599;
assign addr[35708]= 959229189;
assign addr[35709]= 890198924;
assign addr[35710]= 820039373;
assign addr[35711]= 748839539;
assign addr[35712]= 676689746;
assign addr[35713]= 603681519;
assign addr[35714]= 529907477;
assign addr[35715]= 455461206;
assign addr[35716]= 380437148;
assign addr[35717]= 304930476;
assign addr[35718]= 229036977;
assign addr[35719]= 152852926;
assign addr[35720]= 76474970;
assign addr[35721]= 0;
assign addr[35722]= -76474970;
assign addr[35723]= -152852926;
assign addr[35724]= -229036977;
assign addr[35725]= -304930476;
assign addr[35726]= -380437148;
assign addr[35727]= -455461206;
assign addr[35728]= -529907477;
assign addr[35729]= -603681519;
assign addr[35730]= -676689746;
assign addr[35731]= -748839539;
assign addr[35732]= -820039373;
assign addr[35733]= -890198924;
assign addr[35734]= -959229189;
assign addr[35735]= -1027042599;
assign addr[35736]= -1093553126;
assign addr[35737]= -1158676398;
assign addr[35738]= -1222329801;
assign addr[35739]= -1284432584;
assign addr[35740]= -1344905966;
assign addr[35741]= -1403673233;
assign addr[35742]= -1460659832;
assign addr[35743]= -1515793473;
assign addr[35744]= -1569004214;
assign addr[35745]= -1620224553;
assign addr[35746]= -1669389513;
assign addr[35747]= -1716436725;
assign addr[35748]= -1761306505;
assign addr[35749]= -1803941934;
assign addr[35750]= -1844288924;
assign addr[35751]= -1882296293;
assign addr[35752]= -1917915825;
assign addr[35753]= -1951102334;
assign addr[35754]= -1981813720;
assign addr[35755]= -2010011024;
assign addr[35756]= -2035658475;
assign addr[35757]= -2058723538;
assign addr[35758]= -2079176953;
assign addr[35759]= -2096992772;
assign addr[35760]= -2112148396;
assign addr[35761]= -2124624598;
assign addr[35762]= -2134405552;
assign addr[35763]= -2141478848;
assign addr[35764]= -2145835515;
assign addr[35765]= -2147470025;
assign addr[35766]= -2146380306;
assign addr[35767]= -2142567738;
assign addr[35768]= -2136037160;
assign addr[35769]= -2126796855;
assign addr[35770]= -2114858546;
assign addr[35771]= -2100237377;
assign addr[35772]= -2082951896;
assign addr[35773]= -2063024031;
assign addr[35774]= -2040479063;
assign addr[35775]= -2015345591;
assign addr[35776]= -1987655498;
assign addr[35777]= -1957443913;
assign addr[35778]= -1924749160;
assign addr[35779]= -1889612716;
assign addr[35780]= -1852079154;
assign addr[35781]= -1812196087;
assign addr[35782]= -1770014111;
assign addr[35783]= -1725586737;
assign addr[35784]= -1678970324;
assign addr[35785]= -1630224009;
assign addr[35786]= -1579409630;
assign addr[35787]= -1526591649;
assign addr[35788]= -1471837070;
assign addr[35789]= -1415215352;
assign addr[35790]= -1356798326;
assign addr[35791]= -1296660098;
assign addr[35792]= -1234876957;
assign addr[35793]= -1171527280;
assign addr[35794]= -1106691431;
assign addr[35795]= -1040451659;
assign addr[35796]= -972891995;
assign addr[35797]= -904098143;
assign addr[35798]= -834157373;
assign addr[35799]= -763158411;
assign addr[35800]= -691191324;
assign addr[35801]= -618347408;
assign addr[35802]= -544719071;
assign addr[35803]= -470399716;
assign addr[35804]= -395483624;
assign addr[35805]= -320065829;
assign addr[35806]= -244242007;
assign addr[35807]= -168108346;
assign addr[35808]= -91761426;
assign addr[35809]= -15298099;
assign addr[35810]= 61184634;
assign addr[35811]= 137589750;
assign addr[35812]= 213820322;
assign addr[35813]= 289779648;
assign addr[35814]= 365371365;
assign addr[35815]= 440499581;
assign addr[35816]= 515068990;
assign addr[35817]= 588984994;
assign addr[35818]= 662153826;
assign addr[35819]= 734482665;
assign addr[35820]= 805879757;
assign addr[35821]= 876254528;
assign addr[35822]= 945517704;
assign addr[35823]= 1013581418;
assign addr[35824]= 1080359326;
assign addr[35825]= 1145766716;
assign addr[35826]= 1209720613;
assign addr[35827]= 1272139887;
assign addr[35828]= 1332945355;
assign addr[35829]= 1392059879;
assign addr[35830]= 1449408469;
assign addr[35831]= 1504918373;
assign addr[35832]= 1558519173;
assign addr[35833]= 1610142873;
assign addr[35834]= 1659723983;
assign addr[35835]= 1707199606;
assign addr[35836]= 1752509516;
assign addr[35837]= 1795596234;
assign addr[35838]= 1836405100;
assign addr[35839]= 1874884346;
assign addr[35840]= 1910985158;
assign addr[35841]= 1944661739;
assign addr[35842]= 1975871368;
assign addr[35843]= 2004574453;
assign addr[35844]= 2030734582;
assign addr[35845]= 2054318569;
assign addr[35846]= 2075296495;
assign addr[35847]= 2093641749;
assign addr[35848]= 2109331059;
assign addr[35849]= 2122344521;
assign addr[35850]= 2132665626;
assign addr[35851]= 2140281282;
assign addr[35852]= 2145181827;
assign addr[35853]= 2147361045;
assign addr[35854]= 2146816171;
assign addr[35855]= 2143547897;
assign addr[35856]= 2137560369;
assign addr[35857]= 2128861181;
assign addr[35858]= 2117461370;
assign addr[35859]= 2103375398;
assign addr[35860]= 2086621133;
assign addr[35861]= 2067219829;
assign addr[35862]= 2045196100;
assign addr[35863]= 2020577882;
assign addr[35864]= 1993396407;
assign addr[35865]= 1963686155;
assign addr[35866]= 1931484818;
assign addr[35867]= 1896833245;
assign addr[35868]= 1859775393;
assign addr[35869]= 1820358275;
assign addr[35870]= 1778631892;
assign addr[35871]= 1734649179;
assign addr[35872]= 1688465931;
assign addr[35873]= 1640140734;
assign addr[35874]= 1589734894;
assign addr[35875]= 1537312353;
assign addr[35876]= 1482939614;
assign addr[35877]= 1426685652;
assign addr[35878]= 1368621831;
assign addr[35879]= 1308821808;
assign addr[35880]= 1247361445;
assign addr[35881]= 1184318708;
assign addr[35882]= 1119773573;
assign addr[35883]= 1053807919;
assign addr[35884]= 986505429;
assign addr[35885]= 917951481;
assign addr[35886]= 848233042;
assign addr[35887]= 777438554;
assign addr[35888]= 705657826;
assign addr[35889]= 632981917;
assign addr[35890]= 559503022;
assign addr[35891]= 485314355;
assign addr[35892]= 410510029;
assign addr[35893]= 335184940;
assign addr[35894]= 259434643;
assign addr[35895]= 183355234;
assign addr[35896]= 107043224;
assign addr[35897]= 30595422;
assign addr[35898]= -45891193;
assign addr[35899]= -122319591;
assign addr[35900]= -198592817;
assign addr[35901]= -274614114;
assign addr[35902]= -350287041;
assign addr[35903]= -425515602;
assign addr[35904]= -500204365;
assign addr[35905]= -574258580;
assign addr[35906]= -647584304;
assign addr[35907]= -720088517;
assign addr[35908]= -791679244;
assign addr[35909]= -862265664;
assign addr[35910]= -931758235;
assign addr[35911]= -1000068799;
assign addr[35912]= -1067110699;
assign addr[35913]= -1132798888;
assign addr[35914]= -1197050035;
assign addr[35915]= -1259782632;
assign addr[35916]= -1320917099;
assign addr[35917]= -1380375881;
assign addr[35918]= -1438083551;
assign addr[35919]= -1493966902;
assign addr[35920]= -1547955041;
assign addr[35921]= -1599979481;
assign addr[35922]= -1649974225;
assign addr[35923]= -1697875851;
assign addr[35924]= -1743623590;
assign addr[35925]= -1787159411;
assign addr[35926]= -1828428082;
assign addr[35927]= -1867377253;
assign addr[35928]= -1903957513;
assign addr[35929]= -1938122457;
assign addr[35930]= -1969828744;
assign addr[35931]= -1999036154;
assign addr[35932]= -2025707632;
assign addr[35933]= -2049809346;
assign addr[35934]= -2071310720;
assign addr[35935]= -2090184478;
assign addr[35936]= -2106406677;
assign addr[35937]= -2119956737;
assign addr[35938]= -2130817471;
assign addr[35939]= -2138975100;
assign addr[35940]= -2144419275;
assign addr[35941]= -2147143090;
assign addr[35942]= -2147143090;
assign addr[35943]= -2144419275;
assign addr[35944]= -2138975100;
assign addr[35945]= -2130817471;
assign addr[35946]= -2119956737;
assign addr[35947]= -2106406677;
assign addr[35948]= -2090184478;
assign addr[35949]= -2071310720;
assign addr[35950]= -2049809346;
assign addr[35951]= -2025707632;
assign addr[35952]= -1999036154;
assign addr[35953]= -1969828744;
assign addr[35954]= -1938122457;
assign addr[35955]= -1903957513;
assign addr[35956]= -1867377253;
assign addr[35957]= -1828428082;
assign addr[35958]= -1787159411;
assign addr[35959]= -1743623590;
assign addr[35960]= -1697875851;
assign addr[35961]= -1649974225;
assign addr[35962]= -1599979481;
assign addr[35963]= -1547955041;
assign addr[35964]= -1493966902;
assign addr[35965]= -1438083551;
assign addr[35966]= -1380375881;
assign addr[35967]= -1320917099;
assign addr[35968]= -1259782632;
assign addr[35969]= -1197050035;
assign addr[35970]= -1132798888;
assign addr[35971]= -1067110699;
assign addr[35972]= -1000068799;
assign addr[35973]= -931758235;
assign addr[35974]= -862265664;
assign addr[35975]= -791679244;
assign addr[35976]= -720088517;
assign addr[35977]= -647584304;
assign addr[35978]= -574258580;
assign addr[35979]= -500204365;
assign addr[35980]= -425515602;
assign addr[35981]= -350287041;
assign addr[35982]= -274614114;
assign addr[35983]= -198592817;
assign addr[35984]= -122319591;
assign addr[35985]= -45891193;
assign addr[35986]= 30595422;
assign addr[35987]= 107043224;
assign addr[35988]= 183355234;
assign addr[35989]= 259434643;
assign addr[35990]= 335184940;
assign addr[35991]= 410510029;
assign addr[35992]= 485314355;
assign addr[35993]= 559503022;
assign addr[35994]= 632981917;
assign addr[35995]= 705657826;
assign addr[35996]= 777438554;
assign addr[35997]= 848233042;
assign addr[35998]= 917951481;
assign addr[35999]= 986505429;
assign addr[36000]= 1053807919;
assign addr[36001]= 1119773573;
assign addr[36002]= 1184318708;
assign addr[36003]= 1247361445;
assign addr[36004]= 1308821808;
assign addr[36005]= 1368621831;
assign addr[36006]= 1426685652;
assign addr[36007]= 1482939614;
assign addr[36008]= 1537312353;
assign addr[36009]= 1589734894;
assign addr[36010]= 1640140734;
assign addr[36011]= 1688465931;
assign addr[36012]= 1734649179;
assign addr[36013]= 1778631892;
assign addr[36014]= 1820358275;
assign addr[36015]= 1859775393;
assign addr[36016]= 1896833245;
assign addr[36017]= 1931484818;
assign addr[36018]= 1963686155;
assign addr[36019]= 1993396407;
assign addr[36020]= 2020577882;
assign addr[36021]= 2045196100;
assign addr[36022]= 2067219829;
assign addr[36023]= 2086621133;
assign addr[36024]= 2103375398;
assign addr[36025]= 2117461370;
assign addr[36026]= 2128861181;
assign addr[36027]= 2137560369;
assign addr[36028]= 2143547897;
assign addr[36029]= 2146816171;
assign addr[36030]= 2147361045;
assign addr[36031]= 2145181827;
assign addr[36032]= 2140281282;
assign addr[36033]= 2132665626;
assign addr[36034]= 2122344521;
assign addr[36035]= 2109331059;
assign addr[36036]= 2093641749;
assign addr[36037]= 2075296495;
assign addr[36038]= 2054318569;
assign addr[36039]= 2030734582;
assign addr[36040]= 2004574453;
assign addr[36041]= 1975871368;
assign addr[36042]= 1944661739;
assign addr[36043]= 1910985158;
assign addr[36044]= 1874884346;
assign addr[36045]= 1836405100;
assign addr[36046]= 1795596234;
assign addr[36047]= 1752509516;
assign addr[36048]= 1707199606;
assign addr[36049]= 1659723983;
assign addr[36050]= 1610142873;
assign addr[36051]= 1558519173;
assign addr[36052]= 1504918373;
assign addr[36053]= 1449408469;
assign addr[36054]= 1392059879;
assign addr[36055]= 1332945355;
assign addr[36056]= 1272139887;
assign addr[36057]= 1209720613;
assign addr[36058]= 1145766716;
assign addr[36059]= 1080359326;
assign addr[36060]= 1013581418;
assign addr[36061]= 945517704;
assign addr[36062]= 876254528;
assign addr[36063]= 805879757;
assign addr[36064]= 734482665;
assign addr[36065]= 662153826;
assign addr[36066]= 588984994;
assign addr[36067]= 515068990;
assign addr[36068]= 440499581;
assign addr[36069]= 365371365;
assign addr[36070]= 289779648;
assign addr[36071]= 213820322;
assign addr[36072]= 137589750;
assign addr[36073]= 61184634;
assign addr[36074]= -15298099;
assign addr[36075]= -91761426;
assign addr[36076]= -168108346;
assign addr[36077]= -244242007;
assign addr[36078]= -320065829;
assign addr[36079]= -395483624;
assign addr[36080]= -470399716;
assign addr[36081]= -544719071;
assign addr[36082]= -618347408;
assign addr[36083]= -691191324;
assign addr[36084]= -763158411;
assign addr[36085]= -834157373;
assign addr[36086]= -904098143;
assign addr[36087]= -972891995;
assign addr[36088]= -1040451659;
assign addr[36089]= -1106691431;
assign addr[36090]= -1171527280;
assign addr[36091]= -1234876957;
assign addr[36092]= -1296660098;
assign addr[36093]= -1356798326;
assign addr[36094]= -1415215352;
assign addr[36095]= -1471837070;
assign addr[36096]= -1526591649;
assign addr[36097]= -1579409630;
assign addr[36098]= -1630224009;
assign addr[36099]= -1678970324;
assign addr[36100]= -1725586737;
assign addr[36101]= -1770014111;
assign addr[36102]= -1812196087;
assign addr[36103]= -1852079154;
assign addr[36104]= -1889612716;
assign addr[36105]= -1924749160;
assign addr[36106]= -1957443913;
assign addr[36107]= -1987655498;
assign addr[36108]= -2015345591;
assign addr[36109]= -2040479063;
assign addr[36110]= -2063024031;
assign addr[36111]= -2082951896;
assign addr[36112]= -2100237377;
assign addr[36113]= -2114858546;
assign addr[36114]= -2126796855;
assign addr[36115]= -2136037160;
assign addr[36116]= -2142567738;
assign addr[36117]= -2146380306;
assign addr[36118]= -2147470025;
assign addr[36119]= -2145835515;
assign addr[36120]= -2141478848;
assign addr[36121]= -2134405552;
assign addr[36122]= -2124624598;
assign addr[36123]= -2112148396;
assign addr[36124]= -2096992772;
assign addr[36125]= -2079176953;
assign addr[36126]= -2058723538;
assign addr[36127]= -2035658475;
assign addr[36128]= -2010011024;
assign addr[36129]= -1981813720;
assign addr[36130]= -1951102334;
assign addr[36131]= -1917915825;
assign addr[36132]= -1882296293;
assign addr[36133]= -1844288924;
assign addr[36134]= -1803941934;
assign addr[36135]= -1761306505;
assign addr[36136]= -1716436725;
assign addr[36137]= -1669389513;
assign addr[36138]= -1620224553;
assign addr[36139]= -1569004214;
assign addr[36140]= -1515793473;
assign addr[36141]= -1460659832;
assign addr[36142]= -1403673233;
assign addr[36143]= -1344905966;
assign addr[36144]= -1284432584;
assign addr[36145]= -1222329801;
assign addr[36146]= -1158676398;
assign addr[36147]= -1093553126;
assign addr[36148]= -1027042599;
assign addr[36149]= -959229189;
assign addr[36150]= -890198924;
assign addr[36151]= -820039373;
assign addr[36152]= -748839539;
assign addr[36153]= -676689746;
assign addr[36154]= -603681519;
assign addr[36155]= -529907477;
assign addr[36156]= -455461206;
assign addr[36157]= -380437148;
assign addr[36158]= -304930476;
assign addr[36159]= -229036977;
assign addr[36160]= -152852926;
assign addr[36161]= -76474970;
assign addr[36162]= 0;
assign addr[36163]= 76474970;
assign addr[36164]= 152852926;
assign addr[36165]= 229036977;
assign addr[36166]= 304930476;
assign addr[36167]= 380437148;
assign addr[36168]= 455461206;
assign addr[36169]= 529907477;
assign addr[36170]= 603681519;
assign addr[36171]= 676689746;
assign addr[36172]= 748839539;
assign addr[36173]= 820039373;
assign addr[36174]= 890198924;
assign addr[36175]= 959229189;
assign addr[36176]= 1027042599;
assign addr[36177]= 1093553126;
assign addr[36178]= 1158676398;
assign addr[36179]= 1222329801;
assign addr[36180]= 1284432584;
assign addr[36181]= 1344905966;
assign addr[36182]= 1403673233;
assign addr[36183]= 1460659832;
assign addr[36184]= 1515793473;
assign addr[36185]= 1569004214;
assign addr[36186]= 1620224553;
assign addr[36187]= 1669389513;
assign addr[36188]= 1716436725;
assign addr[36189]= 1761306505;
assign addr[36190]= 1803941934;
assign addr[36191]= 1844288924;
assign addr[36192]= 1882296293;
assign addr[36193]= 1917915825;
assign addr[36194]= 1951102334;
assign addr[36195]= 1981813720;
assign addr[36196]= 2010011024;
assign addr[36197]= 2035658475;
assign addr[36198]= 2058723538;
assign addr[36199]= 2079176953;
assign addr[36200]= 2096992772;
assign addr[36201]= 2112148396;
assign addr[36202]= 2124624598;
assign addr[36203]= 2134405552;
assign addr[36204]= 2141478848;
assign addr[36205]= 2145835515;
assign addr[36206]= 2147470025;
assign addr[36207]= 2146380306;
assign addr[36208]= 2142567738;
assign addr[36209]= 2136037160;
assign addr[36210]= 2126796855;
assign addr[36211]= 2114858546;
assign addr[36212]= 2100237377;
assign addr[36213]= 2082951896;
assign addr[36214]= 2063024031;
assign addr[36215]= 2040479063;
assign addr[36216]= 2015345591;
assign addr[36217]= 1987655498;
assign addr[36218]= 1957443913;
assign addr[36219]= 1924749160;
assign addr[36220]= 1889612716;
assign addr[36221]= 1852079154;
assign addr[36222]= 1812196087;
assign addr[36223]= 1770014111;
assign addr[36224]= 1725586737;
assign addr[36225]= 1678970324;
assign addr[36226]= 1630224009;
assign addr[36227]= 1579409630;
assign addr[36228]= 1526591649;
assign addr[36229]= 1471837070;
assign addr[36230]= 1415215352;
assign addr[36231]= 1356798326;
assign addr[36232]= 1296660098;
assign addr[36233]= 1234876957;
assign addr[36234]= 1171527280;
assign addr[36235]= 1106691431;
assign addr[36236]= 1040451659;
assign addr[36237]= 972891995;
assign addr[36238]= 904098143;
assign addr[36239]= 834157373;
assign addr[36240]= 763158411;
assign addr[36241]= 691191324;
assign addr[36242]= 618347408;
assign addr[36243]= 544719071;
assign addr[36244]= 470399716;
assign addr[36245]= 395483624;
assign addr[36246]= 320065829;
assign addr[36247]= 244242007;
assign addr[36248]= 168108346;
assign addr[36249]= 91761426;
assign addr[36250]= 15298099;
assign addr[36251]= -61184634;
assign addr[36252]= -137589750;
assign addr[36253]= -213820322;
assign addr[36254]= -289779648;
assign addr[36255]= -365371365;
assign addr[36256]= -440499581;
assign addr[36257]= -515068990;
assign addr[36258]= -588984994;
assign addr[36259]= -662153826;
assign addr[36260]= -734482665;
assign addr[36261]= -805879757;
assign addr[36262]= -876254528;
assign addr[36263]= -945517704;
assign addr[36264]= -1013581418;
assign addr[36265]= -1080359326;
assign addr[36266]= -1145766716;
assign addr[36267]= -1209720613;
assign addr[36268]= -1272139887;
assign addr[36269]= -1332945355;
assign addr[36270]= -1392059879;
assign addr[36271]= -1449408469;
assign addr[36272]= -1504918373;
assign addr[36273]= -1558519173;
assign addr[36274]= -1610142873;
assign addr[36275]= -1659723983;
assign addr[36276]= -1707199606;
assign addr[36277]= -1752509516;
assign addr[36278]= -1795596234;
assign addr[36279]= -1836405100;
assign addr[36280]= -1874884346;
assign addr[36281]= -1910985158;
assign addr[36282]= -1944661739;
assign addr[36283]= -1975871368;
assign addr[36284]= -2004574453;
assign addr[36285]= -2030734582;
assign addr[36286]= -2054318569;
assign addr[36287]= -2075296495;
assign addr[36288]= -2093641749;
assign addr[36289]= -2109331059;
assign addr[36290]= -2122344521;
assign addr[36291]= -2132665626;
assign addr[36292]= -2140281282;
assign addr[36293]= -2145181827;
assign addr[36294]= -2147361045;
assign addr[36295]= -2146816171;
assign addr[36296]= -2143547897;
assign addr[36297]= -2137560369;
assign addr[36298]= -2128861181;
assign addr[36299]= -2117461370;
assign addr[36300]= -2103375398;
assign addr[36301]= -2086621133;
assign addr[36302]= -2067219829;
assign addr[36303]= -2045196100;
assign addr[36304]= -2020577882;
assign addr[36305]= -1993396407;
assign addr[36306]= -1963686155;
assign addr[36307]= -1931484818;
assign addr[36308]= -1896833245;
assign addr[36309]= -1859775393;
assign addr[36310]= -1820358275;
assign addr[36311]= -1778631892;
assign addr[36312]= -1734649179;
assign addr[36313]= -1688465931;
assign addr[36314]= -1640140734;
assign addr[36315]= -1589734894;
assign addr[36316]= -1537312353;
assign addr[36317]= -1482939614;
assign addr[36318]= -1426685652;
assign addr[36319]= -1368621831;
assign addr[36320]= -1308821808;
assign addr[36321]= -1247361445;
assign addr[36322]= -1184318708;
assign addr[36323]= -1119773573;
assign addr[36324]= -1053807919;
assign addr[36325]= -986505429;
assign addr[36326]= -917951481;
assign addr[36327]= -848233042;
assign addr[36328]= -777438554;
assign addr[36329]= -705657826;
assign addr[36330]= -632981917;
assign addr[36331]= -559503022;
assign addr[36332]= -485314355;
assign addr[36333]= -410510029;
assign addr[36334]= -335184940;
assign addr[36335]= -259434643;
assign addr[36336]= -183355234;
assign addr[36337]= -107043224;
assign addr[36338]= -30595422;
assign addr[36339]= 45891193;
assign addr[36340]= 122319591;
assign addr[36341]= 198592817;
assign addr[36342]= 274614114;
assign addr[36343]= 350287041;
assign addr[36344]= 425515602;
assign addr[36345]= 500204365;
assign addr[36346]= 574258580;
assign addr[36347]= 647584304;
assign addr[36348]= 720088517;
assign addr[36349]= 791679244;
assign addr[36350]= 862265664;
assign addr[36351]= 931758235;
assign addr[36352]= 1000068799;
assign addr[36353]= 1067110699;
assign addr[36354]= 1132798888;
assign addr[36355]= 1197050035;
assign addr[36356]= 1259782632;
assign addr[36357]= 1320917099;
assign addr[36358]= 1380375881;
assign addr[36359]= 1438083551;
assign addr[36360]= 1493966902;
assign addr[36361]= 1547955041;
assign addr[36362]= 1599979481;
assign addr[36363]= 1649974225;
assign addr[36364]= 1697875851;
assign addr[36365]= 1743623590;
assign addr[36366]= 1787159411;
assign addr[36367]= 1828428082;
assign addr[36368]= 1867377253;
assign addr[36369]= 1903957513;
assign addr[36370]= 1938122457;
assign addr[36371]= 1969828744;
assign addr[36372]= 1999036154;
assign addr[36373]= 2025707632;
assign addr[36374]= 2049809346;
assign addr[36375]= 2071310720;
assign addr[36376]= 2090184478;
assign addr[36377]= 2106406677;
assign addr[36378]= 2119956737;
assign addr[36379]= 2130817471;
assign addr[36380]= 2138975100;
assign addr[36381]= 2144419275;
assign addr[36382]= 2147143090;
assign addr[36383]= 2147143090;
assign addr[36384]= 2144419275;
assign addr[36385]= 2138975100;
assign addr[36386]= 2130817471;
assign addr[36387]= 2119956737;
assign addr[36388]= 2106406677;
assign addr[36389]= 2090184478;
assign addr[36390]= 2071310720;
assign addr[36391]= 2049809346;
assign addr[36392]= 2025707632;
assign addr[36393]= 1999036154;
assign addr[36394]= 1969828744;
assign addr[36395]= 1938122457;
assign addr[36396]= 1903957513;
assign addr[36397]= 1867377253;
assign addr[36398]= 1828428082;
assign addr[36399]= 1787159411;
assign addr[36400]= 1743623590;
assign addr[36401]= 1697875851;
assign addr[36402]= 1649974225;
assign addr[36403]= 1599979481;
assign addr[36404]= 1547955041;
assign addr[36405]= 1493966902;
assign addr[36406]= 1438083551;
assign addr[36407]= 1380375881;
assign addr[36408]= 1320917099;
assign addr[36409]= 1259782632;
assign addr[36410]= 1197050035;
assign addr[36411]= 1132798888;
assign addr[36412]= 1067110699;
assign addr[36413]= 1000068799;
assign addr[36414]= 931758235;
assign addr[36415]= 862265664;
assign addr[36416]= 791679244;
assign addr[36417]= 720088517;
assign addr[36418]= 647584304;
assign addr[36419]= 574258580;
assign addr[36420]= 500204365;
assign addr[36421]= 425515602;
assign addr[36422]= 350287041;
assign addr[36423]= 274614114;
assign addr[36424]= 198592817;
assign addr[36425]= 122319591;
assign addr[36426]= 45891193;
assign addr[36427]= -30595422;
assign addr[36428]= -107043224;
assign addr[36429]= -183355234;
assign addr[36430]= -259434643;
assign addr[36431]= -335184940;
assign addr[36432]= -410510029;
assign addr[36433]= -485314355;
assign addr[36434]= -559503022;
assign addr[36435]= -632981917;
assign addr[36436]= -705657826;
assign addr[36437]= -777438554;
assign addr[36438]= -848233042;
assign addr[36439]= -917951481;
assign addr[36440]= -986505429;
assign addr[36441]= -1053807919;
assign addr[36442]= -1119773573;
assign addr[36443]= -1184318708;
assign addr[36444]= -1247361445;
assign addr[36445]= -1308821808;
assign addr[36446]= -1368621831;
assign addr[36447]= -1426685652;
assign addr[36448]= -1482939614;
assign addr[36449]= -1537312353;
assign addr[36450]= -1589734894;
assign addr[36451]= -1640140734;
assign addr[36452]= -1688465931;
assign addr[36453]= -1734649179;
assign addr[36454]= -1778631892;
assign addr[36455]= -1820358275;
assign addr[36456]= -1859775393;
assign addr[36457]= -1896833245;
assign addr[36458]= -1931484818;
assign addr[36459]= -1963686155;
assign addr[36460]= -1993396407;
assign addr[36461]= -2020577882;
assign addr[36462]= -2045196100;
assign addr[36463]= -2067219829;
assign addr[36464]= -2086621133;
assign addr[36465]= -2103375398;
assign addr[36466]= -2117461370;
assign addr[36467]= -2128861181;
assign addr[36468]= -2137560369;
assign addr[36469]= -2143547897;
assign addr[36470]= -2146816171;
assign addr[36471]= -2147361045;
assign addr[36472]= -2145181827;
assign addr[36473]= -2140281282;
assign addr[36474]= -2132665626;
assign addr[36475]= -2122344521;
assign addr[36476]= -2109331059;
assign addr[36477]= -2093641749;
assign addr[36478]= -2075296495;
assign addr[36479]= -2054318569;
assign addr[36480]= -2030734582;
assign addr[36481]= -2004574453;
assign addr[36482]= -1975871368;
assign addr[36483]= -1944661739;
assign addr[36484]= -1910985158;
assign addr[36485]= -1874884346;
assign addr[36486]= -1836405100;
assign addr[36487]= -1795596234;
assign addr[36488]= -1752509516;
assign addr[36489]= -1707199606;
assign addr[36490]= -1659723983;
assign addr[36491]= -1610142873;
assign addr[36492]= -1558519173;
assign addr[36493]= -1504918373;
assign addr[36494]= -1449408469;
assign addr[36495]= -1392059879;
assign addr[36496]= -1332945355;
assign addr[36497]= -1272139887;
assign addr[36498]= -1209720613;
assign addr[36499]= -1145766716;
assign addr[36500]= -1080359326;
assign addr[36501]= -1013581418;
assign addr[36502]= -945517704;
assign addr[36503]= -876254528;
assign addr[36504]= -805879757;
assign addr[36505]= -734482665;
assign addr[36506]= -662153826;
assign addr[36507]= -588984994;
assign addr[36508]= -515068990;
assign addr[36509]= -440499581;
assign addr[36510]= -365371365;
assign addr[36511]= -289779648;
assign addr[36512]= -213820322;
assign addr[36513]= -137589750;
assign addr[36514]= -61184634;
assign addr[36515]= 15298099;
assign addr[36516]= 91761426;
assign addr[36517]= 168108346;
assign addr[36518]= 244242007;
assign addr[36519]= 320065829;
assign addr[36520]= 395483624;
assign addr[36521]= 470399716;
assign addr[36522]= 544719071;
assign addr[36523]= 618347408;
assign addr[36524]= 691191324;
assign addr[36525]= 763158411;
assign addr[36526]= 834157373;
assign addr[36527]= 904098143;
assign addr[36528]= 972891995;
assign addr[36529]= 1040451659;
assign addr[36530]= 1106691431;
assign addr[36531]= 1171527280;
assign addr[36532]= 1234876957;
assign addr[36533]= 1296660098;
assign addr[36534]= 1356798326;
assign addr[36535]= 1415215352;
assign addr[36536]= 1471837070;
assign addr[36537]= 1526591649;
assign addr[36538]= 1579409630;
assign addr[36539]= 1630224009;
assign addr[36540]= 1678970324;
assign addr[36541]= 1725586737;
assign addr[36542]= 1770014111;
assign addr[36543]= 1812196087;
assign addr[36544]= 1852079154;
assign addr[36545]= 1889612716;
assign addr[36546]= 1924749160;
assign addr[36547]= 1957443913;
assign addr[36548]= 1987655498;
assign addr[36549]= 2015345591;
assign addr[36550]= 2040479063;
assign addr[36551]= 2063024031;
assign addr[36552]= 2082951896;
assign addr[36553]= 2100237377;
assign addr[36554]= 2114858546;
assign addr[36555]= 2126796855;
assign addr[36556]= 2136037160;
assign addr[36557]= 2142567738;
assign addr[36558]= 2146380306;
assign addr[36559]= 2147470025;
assign addr[36560]= 2145835515;
assign addr[36561]= 2141478848;
assign addr[36562]= 2134405552;
assign addr[36563]= 2124624598;
assign addr[36564]= 2112148396;
assign addr[36565]= 2096992772;
assign addr[36566]= 2079176953;
assign addr[36567]= 2058723538;
assign addr[36568]= 2035658475;
assign addr[36569]= 2010011024;
assign addr[36570]= 1981813720;
assign addr[36571]= 1951102334;
assign addr[36572]= 1917915825;
assign addr[36573]= 1882296293;
assign addr[36574]= 1844288924;
assign addr[36575]= 1803941934;
assign addr[36576]= 1761306505;
assign addr[36577]= 1716436725;
assign addr[36578]= 1669389513;
assign addr[36579]= 1620224553;
assign addr[36580]= 1569004214;
assign addr[36581]= 1515793473;
assign addr[36582]= 1460659832;
assign addr[36583]= 1403673233;
assign addr[36584]= 1344905966;
assign addr[36585]= 1284432584;
assign addr[36586]= 1222329801;
assign addr[36587]= 1158676398;
assign addr[36588]= 1093553126;
assign addr[36589]= 1027042599;
assign addr[36590]= 959229189;
assign addr[36591]= 890198924;
assign addr[36592]= 820039373;
assign addr[36593]= 748839539;
assign addr[36594]= 676689746;
assign addr[36595]= 603681519;
assign addr[36596]= 529907477;
assign addr[36597]= 455461206;
assign addr[36598]= 380437148;
assign addr[36599]= 304930476;
assign addr[36600]= 229036977;
assign addr[36601]= 152852926;
assign addr[36602]= 76474970;
assign addr[36603]= 0;
assign addr[36604]= -76474970;
assign addr[36605]= -152852926;
assign addr[36606]= -229036977;
assign addr[36607]= -304930476;
assign addr[36608]= -380437148;
assign addr[36609]= -455461206;
assign addr[36610]= -529907477;
assign addr[36611]= -603681519;
assign addr[36612]= -676689746;
assign addr[36613]= -748839539;
assign addr[36614]= -820039373;
assign addr[36615]= -890198924;
assign addr[36616]= -959229189;
assign addr[36617]= -1027042599;
assign addr[36618]= -1093553126;
assign addr[36619]= -1158676398;
assign addr[36620]= -1222329801;
assign addr[36621]= -1284432584;
assign addr[36622]= -1344905966;
assign addr[36623]= -1403673233;
assign addr[36624]= -1460659832;
assign addr[36625]= -1515793473;
assign addr[36626]= -1569004214;
assign addr[36627]= -1620224553;
assign addr[36628]= -1669389513;
assign addr[36629]= -1716436725;
assign addr[36630]= -1761306505;
assign addr[36631]= -1803941934;
assign addr[36632]= -1844288924;
assign addr[36633]= -1882296293;
assign addr[36634]= -1917915825;
assign addr[36635]= -1951102334;
assign addr[36636]= -1981813720;
assign addr[36637]= -2010011024;
assign addr[36638]= -2035658475;
assign addr[36639]= -2058723538;
assign addr[36640]= -2079176953;
assign addr[36641]= -2096992772;
assign addr[36642]= -2112148396;
assign addr[36643]= -2124624598;
assign addr[36644]= -2134405552;
assign addr[36645]= -2141478848;
assign addr[36646]= -2145835515;
assign addr[36647]= -2147470025;
assign addr[36648]= -2146380306;
assign addr[36649]= -2142567738;
assign addr[36650]= -2136037160;
assign addr[36651]= -2126796855;
assign addr[36652]= -2114858546;
assign addr[36653]= -2100237377;
assign addr[36654]= -2082951896;
assign addr[36655]= -2063024031;
assign addr[36656]= -2040479063;
assign addr[36657]= -2015345591;
assign addr[36658]= -1987655498;
assign addr[36659]= -1957443913;
assign addr[36660]= -1924749160;
assign addr[36661]= -1889612716;
assign addr[36662]= -1852079154;
assign addr[36663]= -1812196087;
assign addr[36664]= -1770014111;
assign addr[36665]= -1725586737;
assign addr[36666]= -1678970324;
assign addr[36667]= -1630224009;
assign addr[36668]= -1579409630;
assign addr[36669]= -1526591649;
assign addr[36670]= -1471837070;
assign addr[36671]= -1415215352;
assign addr[36672]= -1356798326;
assign addr[36673]= -1296660098;
assign addr[36674]= -1234876957;
assign addr[36675]= -1171527280;
assign addr[36676]= -1106691431;
assign addr[36677]= -1040451659;
assign addr[36678]= -972891995;
assign addr[36679]= -904098143;
assign addr[36680]= -834157373;
assign addr[36681]= -763158411;
assign addr[36682]= -691191324;
assign addr[36683]= -618347408;
assign addr[36684]= -544719071;
assign addr[36685]= -470399716;
assign addr[36686]= -395483624;
assign addr[36687]= -320065829;
assign addr[36688]= -244242007;
assign addr[36689]= -168108346;
assign addr[36690]= -91761426;
assign addr[36691]= -15298099;
assign addr[36692]= 61184634;
assign addr[36693]= 137589750;
assign addr[36694]= 213820322;
assign addr[36695]= 289779648;
assign addr[36696]= 365371365;
assign addr[36697]= 440499581;
assign addr[36698]= 515068990;
assign addr[36699]= 588984994;
assign addr[36700]= 662153826;
assign addr[36701]= 734482665;
assign addr[36702]= 805879757;
assign addr[36703]= 876254528;
assign addr[36704]= 945517704;
assign addr[36705]= 1013581418;
assign addr[36706]= 1080359326;
assign addr[36707]= 1145766716;
assign addr[36708]= 1209720613;
assign addr[36709]= 1272139887;
assign addr[36710]= 1332945355;
assign addr[36711]= 1392059879;
assign addr[36712]= 1449408469;
assign addr[36713]= 1504918373;
assign addr[36714]= 1558519173;
assign addr[36715]= 1610142873;
assign addr[36716]= 1659723983;
assign addr[36717]= 1707199606;
assign addr[36718]= 1752509516;
assign addr[36719]= 1795596234;
assign addr[36720]= 1836405100;
assign addr[36721]= 1874884346;
assign addr[36722]= 1910985158;
assign addr[36723]= 1944661739;
assign addr[36724]= 1975871368;
assign addr[36725]= 2004574453;
assign addr[36726]= 2030734582;
assign addr[36727]= 2054318569;
assign addr[36728]= 2075296495;
assign addr[36729]= 2093641749;
assign addr[36730]= 2109331059;
assign addr[36731]= 2122344521;
assign addr[36732]= 2132665626;
assign addr[36733]= 2140281282;
assign addr[36734]= 2145181827;
assign addr[36735]= 2147361045;
assign addr[36736]= 2146816171;
assign addr[36737]= 2143547897;
assign addr[36738]= 2137560369;
assign addr[36739]= 2128861181;
assign addr[36740]= 2117461370;
assign addr[36741]= 2103375398;
assign addr[36742]= 2086621133;
assign addr[36743]= 2067219829;
assign addr[36744]= 2045196100;
assign addr[36745]= 2020577882;
assign addr[36746]= 1993396407;
assign addr[36747]= 1963686155;
assign addr[36748]= 1931484818;
assign addr[36749]= 1896833245;
assign addr[36750]= 1859775393;
assign addr[36751]= 1820358275;
assign addr[36752]= 1778631892;
assign addr[36753]= 1734649179;
assign addr[36754]= 1688465931;
assign addr[36755]= 1640140734;
assign addr[36756]= 1589734894;
assign addr[36757]= 1537312353;
assign addr[36758]= 1482939614;
assign addr[36759]= 1426685652;
assign addr[36760]= 1368621831;
assign addr[36761]= 1308821808;
assign addr[36762]= 1247361445;
assign addr[36763]= 1184318708;
assign addr[36764]= 1119773573;
assign addr[36765]= 1053807919;
assign addr[36766]= 986505429;
assign addr[36767]= 917951481;
assign addr[36768]= 848233042;
assign addr[36769]= 777438554;
assign addr[36770]= 705657826;
assign addr[36771]= 632981917;
assign addr[36772]= 559503022;
assign addr[36773]= 485314355;
assign addr[36774]= 410510029;
assign addr[36775]= 335184940;
assign addr[36776]= 259434643;
assign addr[36777]= 183355234;
assign addr[36778]= 107043224;
assign addr[36779]= 30595422;
assign addr[36780]= -45891193;
assign addr[36781]= -122319591;
assign addr[36782]= -198592817;
assign addr[36783]= -274614114;
assign addr[36784]= -350287041;
assign addr[36785]= -425515602;
assign addr[36786]= -500204365;
assign addr[36787]= -574258580;
assign addr[36788]= -647584304;
assign addr[36789]= -720088517;
assign addr[36790]= -791679244;
assign addr[36791]= -862265664;
assign addr[36792]= -931758235;
assign addr[36793]= -1000068799;
assign addr[36794]= -1067110699;
assign addr[36795]= -1132798888;
assign addr[36796]= -1197050035;
assign addr[36797]= -1259782632;
assign addr[36798]= -1320917099;
assign addr[36799]= -1380375881;
assign addr[36800]= -1438083551;
assign addr[36801]= -1493966902;
assign addr[36802]= -1547955041;
assign addr[36803]= -1599979481;
assign addr[36804]= -1649974225;
assign addr[36805]= -1697875851;
assign addr[36806]= -1743623590;
assign addr[36807]= -1787159411;
assign addr[36808]= -1828428082;
assign addr[36809]= -1867377253;
assign addr[36810]= -1903957513;
assign addr[36811]= -1938122457;
assign addr[36812]= -1969828744;
assign addr[36813]= -1999036154;
assign addr[36814]= -2025707632;
assign addr[36815]= -2049809346;
assign addr[36816]= -2071310720;
assign addr[36817]= -2090184478;
assign addr[36818]= -2106406677;
assign addr[36819]= -2119956737;
assign addr[36820]= -2130817471;
assign addr[36821]= -2138975100;
assign addr[36822]= -2144419275;
assign addr[36823]= -2147143090;
assign addr[36824]= -2147143090;
assign addr[36825]= -2144419275;
assign addr[36826]= -2138975100;
assign addr[36827]= -2130817471;
assign addr[36828]= -2119956737;
assign addr[36829]= -2106406677;
assign addr[36830]= -2090184478;
assign addr[36831]= -2071310720;
assign addr[36832]= -2049809346;
assign addr[36833]= -2025707632;
assign addr[36834]= -1999036154;
assign addr[36835]= -1969828744;
assign addr[36836]= -1938122457;
assign addr[36837]= -1903957513;
assign addr[36838]= -1867377253;
assign addr[36839]= -1828428082;
assign addr[36840]= -1787159411;
assign addr[36841]= -1743623590;
assign addr[36842]= -1697875851;
assign addr[36843]= -1649974225;
assign addr[36844]= -1599979481;
assign addr[36845]= -1547955041;
assign addr[36846]= -1493966902;
assign addr[36847]= -1438083551;
assign addr[36848]= -1380375881;
assign addr[36849]= -1320917099;
assign addr[36850]= -1259782632;
assign addr[36851]= -1197050035;
assign addr[36852]= -1132798888;
assign addr[36853]= -1067110699;
assign addr[36854]= -1000068799;
assign addr[36855]= -931758235;
assign addr[36856]= -862265664;
assign addr[36857]= -791679244;
assign addr[36858]= -720088517;
assign addr[36859]= -647584304;
assign addr[36860]= -574258580;
assign addr[36861]= -500204365;
assign addr[36862]= -425515602;
assign addr[36863]= -350287041;
assign addr[36864]= -274614114;
assign addr[36865]= -198592817;
assign addr[36866]= -122319591;
assign addr[36867]= -45891193;
assign addr[36868]= 30595422;
assign addr[36869]= 107043224;
assign addr[36870]= 183355234;
assign addr[36871]= 259434643;
assign addr[36872]= 335184940;
assign addr[36873]= 410510029;
assign addr[36874]= 485314355;
assign addr[36875]= 559503022;
assign addr[36876]= 632981917;
assign addr[36877]= 705657826;
assign addr[36878]= 777438554;
assign addr[36879]= 848233042;
assign addr[36880]= 917951481;
assign addr[36881]= 986505429;
assign addr[36882]= 1053807919;
assign addr[36883]= 1119773573;
assign addr[36884]= 1184318708;
assign addr[36885]= 1247361445;
assign addr[36886]= 1308821808;
assign addr[36887]= 1368621831;
assign addr[36888]= 1426685652;
assign addr[36889]= 1482939614;
assign addr[36890]= 1537312353;
assign addr[36891]= 1589734894;
assign addr[36892]= 1640140734;
assign addr[36893]= 1688465931;
assign addr[36894]= 1734649179;
assign addr[36895]= 1778631892;
assign addr[36896]= 1820358275;
assign addr[36897]= 1859775393;
assign addr[36898]= 1896833245;
assign addr[36899]= 1931484818;
assign addr[36900]= 1963686155;
assign addr[36901]= 1993396407;
assign addr[36902]= 2020577882;
assign addr[36903]= 2045196100;
assign addr[36904]= 2067219829;
assign addr[36905]= 2086621133;
assign addr[36906]= 2103375398;
assign addr[36907]= 2117461370;
assign addr[36908]= 2128861181;
assign addr[36909]= 2137560369;
assign addr[36910]= 2143547897;
assign addr[36911]= 2146816171;
assign addr[36912]= 2147361045;
assign addr[36913]= 2145181827;
assign addr[36914]= 2140281282;
assign addr[36915]= 2132665626;
assign addr[36916]= 2122344521;
assign addr[36917]= 2109331059;
assign addr[36918]= 2093641749;
assign addr[36919]= 2075296495;
assign addr[36920]= 2054318569;
assign addr[36921]= 2030734582;
assign addr[36922]= 2004574453;
assign addr[36923]= 1975871368;
assign addr[36924]= 1944661739;
assign addr[36925]= 1910985158;
assign addr[36926]= 1874884346;
assign addr[36927]= 1836405100;
assign addr[36928]= 1795596234;
assign addr[36929]= 1752509516;
assign addr[36930]= 1707199606;
assign addr[36931]= 1659723983;
assign addr[36932]= 1610142873;
assign addr[36933]= 1558519173;
assign addr[36934]= 1504918373;
assign addr[36935]= 1449408469;
assign addr[36936]= 1392059879;
assign addr[36937]= 1332945355;
assign addr[36938]= 1272139887;
assign addr[36939]= 1209720613;
assign addr[36940]= 1145766716;
assign addr[36941]= 1080359326;
assign addr[36942]= 1013581418;
assign addr[36943]= 945517704;
assign addr[36944]= 876254528;
assign addr[36945]= 805879757;
assign addr[36946]= 734482665;
assign addr[36947]= 662153826;
assign addr[36948]= 588984994;
assign addr[36949]= 515068990;
assign addr[36950]= 440499581;
assign addr[36951]= 365371365;
assign addr[36952]= 289779648;
assign addr[36953]= 213820322;
assign addr[36954]= 137589750;
assign addr[36955]= 61184634;
assign addr[36956]= -15298099;
assign addr[36957]= -91761426;
assign addr[36958]= -168108346;
assign addr[36959]= -244242007;
assign addr[36960]= -320065829;
assign addr[36961]= -395483624;
assign addr[36962]= -470399716;
assign addr[36963]= -544719071;
assign addr[36964]= -618347408;
assign addr[36965]= -691191324;
assign addr[36966]= -763158411;
assign addr[36967]= -834157373;
assign addr[36968]= -904098143;
assign addr[36969]= -972891995;
assign addr[36970]= -1040451659;
assign addr[36971]= -1106691431;
assign addr[36972]= -1171527280;
assign addr[36973]= -1234876957;
assign addr[36974]= -1296660098;
assign addr[36975]= -1356798326;
assign addr[36976]= -1415215352;
assign addr[36977]= -1471837070;
assign addr[36978]= -1526591649;
assign addr[36979]= -1579409630;
assign addr[36980]= -1630224009;
assign addr[36981]= -1678970324;
assign addr[36982]= -1725586737;
assign addr[36983]= -1770014111;
assign addr[36984]= -1812196087;
assign addr[36985]= -1852079154;
assign addr[36986]= -1889612716;
assign addr[36987]= -1924749160;
assign addr[36988]= -1957443913;
assign addr[36989]= -1987655498;
assign addr[36990]= -2015345591;
assign addr[36991]= -2040479063;
assign addr[36992]= -2063024031;
assign addr[36993]= -2082951896;
assign addr[36994]= -2100237377;
assign addr[36995]= -2114858546;
assign addr[36996]= -2126796855;
assign addr[36997]= -2136037160;
assign addr[36998]= -2142567738;
assign addr[36999]= -2146380306;
assign addr[37000]= -2147470025;
assign addr[37001]= -2145835515;
assign addr[37002]= -2141478848;
assign addr[37003]= -2134405552;
assign addr[37004]= -2124624598;
assign addr[37005]= -2112148396;
assign addr[37006]= -2096992772;
assign addr[37007]= -2079176953;
assign addr[37008]= -2058723538;
assign addr[37009]= -2035658475;
assign addr[37010]= -2010011024;
assign addr[37011]= -1981813720;
assign addr[37012]= -1951102334;
assign addr[37013]= -1917915825;
assign addr[37014]= -1882296293;
assign addr[37015]= -1844288924;
assign addr[37016]= -1803941934;
assign addr[37017]= -1761306505;
assign addr[37018]= -1716436725;
assign addr[37019]= -1669389513;
assign addr[37020]= -1620224553;
assign addr[37021]= -1569004214;
assign addr[37022]= -1515793473;
assign addr[37023]= -1460659832;
assign addr[37024]= -1403673233;
assign addr[37025]= -1344905966;
assign addr[37026]= -1284432584;
assign addr[37027]= -1222329801;
assign addr[37028]= -1158676398;
assign addr[37029]= -1093553126;
assign addr[37030]= -1027042599;
assign addr[37031]= -959229189;
assign addr[37032]= -890198924;
assign addr[37033]= -820039373;
assign addr[37034]= -748839539;
assign addr[37035]= -676689746;
assign addr[37036]= -603681519;
assign addr[37037]= -529907477;
assign addr[37038]= -455461206;
assign addr[37039]= -380437148;
assign addr[37040]= -304930476;
assign addr[37041]= -229036977;
assign addr[37042]= -152852926;
assign addr[37043]= -76474970;
assign addr[37044]= 0;
assign addr[37045]= 76474970;
assign addr[37046]= 152852926;
assign addr[37047]= 229036977;
assign addr[37048]= 304930476;
assign addr[37049]= 380437148;
assign addr[37050]= 455461206;
assign addr[37051]= 529907477;
assign addr[37052]= 603681519;
assign addr[37053]= 676689746;
assign addr[37054]= 748839539;
assign addr[37055]= 820039373;
assign addr[37056]= 890198924;
assign addr[37057]= 959229189;
assign addr[37058]= 1027042599;
assign addr[37059]= 1093553126;
assign addr[37060]= 1158676398;
assign addr[37061]= 1222329801;
assign addr[37062]= 1284432584;
assign addr[37063]= 1344905966;
assign addr[37064]= 1403673233;
assign addr[37065]= 1460659832;
assign addr[37066]= 1515793473;
assign addr[37067]= 1569004214;
assign addr[37068]= 1620224553;
assign addr[37069]= 1669389513;
assign addr[37070]= 1716436725;
assign addr[37071]= 1761306505;
assign addr[37072]= 1803941934;
assign addr[37073]= 1844288924;
assign addr[37074]= 1882296293;
assign addr[37075]= 1917915825;
assign addr[37076]= 1951102334;
assign addr[37077]= 1981813720;
assign addr[37078]= 2010011024;
assign addr[37079]= 2035658475;
assign addr[37080]= 2058723538;
assign addr[37081]= 2079176953;
assign addr[37082]= 2096992772;
assign addr[37083]= 2112148396;
assign addr[37084]= 2124624598;
assign addr[37085]= 2134405552;
assign addr[37086]= 2141478848;
assign addr[37087]= 2145835515;
assign addr[37088]= 2147470025;
assign addr[37089]= 2146380306;
assign addr[37090]= 2142567738;
assign addr[37091]= 2136037160;
assign addr[37092]= 2126796855;
assign addr[37093]= 2114858546;
assign addr[37094]= 2100237377;
assign addr[37095]= 2082951896;
assign addr[37096]= 2063024031;
assign addr[37097]= 2040479063;
assign addr[37098]= 2015345591;
assign addr[37099]= 1987655498;
assign addr[37100]= 1957443913;
assign addr[37101]= 1924749160;
assign addr[37102]= 1889612716;
assign addr[37103]= 1852079154;
assign addr[37104]= 1812196087;
assign addr[37105]= 1770014111;
assign addr[37106]= 1725586737;
assign addr[37107]= 1678970324;
assign addr[37108]= 1630224009;
assign addr[37109]= 1579409630;
assign addr[37110]= 1526591649;
assign addr[37111]= 1471837070;
assign addr[37112]= 1415215352;
assign addr[37113]= 1356798326;
assign addr[37114]= 1296660098;
assign addr[37115]= 1234876957;
assign addr[37116]= 1171527280;
assign addr[37117]= 1106691431;
assign addr[37118]= 1040451659;
assign addr[37119]= 972891995;
assign addr[37120]= 904098143;
assign addr[37121]= 834157373;
assign addr[37122]= 763158411;
assign addr[37123]= 691191324;
assign addr[37124]= 618347408;
assign addr[37125]= 544719071;
assign addr[37126]= 470399716;
assign addr[37127]= 395483624;
assign addr[37128]= 320065829;
assign addr[37129]= 244242007;
assign addr[37130]= 168108346;
assign addr[37131]= 91761426;
assign addr[37132]= 15298099;
assign addr[37133]= -61184634;
assign addr[37134]= -137589750;
assign addr[37135]= -213820322;
assign addr[37136]= -289779648;
assign addr[37137]= -365371365;
assign addr[37138]= -440499581;
assign addr[37139]= -515068990;
assign addr[37140]= -588984994;
assign addr[37141]= -662153826;
assign addr[37142]= -734482665;
assign addr[37143]= -805879757;
assign addr[37144]= -876254528;
assign addr[37145]= -945517704;
assign addr[37146]= -1013581418;
assign addr[37147]= -1080359326;
assign addr[37148]= -1145766716;
assign addr[37149]= -1209720613;
assign addr[37150]= -1272139887;
assign addr[37151]= -1332945355;
assign addr[37152]= -1392059879;
assign addr[37153]= -1449408469;
assign addr[37154]= -1504918373;
assign addr[37155]= -1558519173;
assign addr[37156]= -1610142873;
assign addr[37157]= -1659723983;
assign addr[37158]= -1707199606;
assign addr[37159]= -1752509516;
assign addr[37160]= -1795596234;
assign addr[37161]= -1836405100;
assign addr[37162]= -1874884346;
assign addr[37163]= -1910985158;
assign addr[37164]= -1944661739;
assign addr[37165]= -1975871368;
assign addr[37166]= -2004574453;
assign addr[37167]= -2030734582;
assign addr[37168]= -2054318569;
assign addr[37169]= -2075296495;
assign addr[37170]= -2093641749;
assign addr[37171]= -2109331059;
assign addr[37172]= -2122344521;
assign addr[37173]= -2132665626;
assign addr[37174]= -2140281282;
assign addr[37175]= -2145181827;
assign addr[37176]= -2147361045;
assign addr[37177]= -2146816171;
assign addr[37178]= -2143547897;
assign addr[37179]= -2137560369;
assign addr[37180]= -2128861181;
assign addr[37181]= -2117461370;
assign addr[37182]= -2103375398;
assign addr[37183]= -2086621133;
assign addr[37184]= -2067219829;
assign addr[37185]= -2045196100;
assign addr[37186]= -2020577882;
assign addr[37187]= -1993396407;
assign addr[37188]= -1963686155;
assign addr[37189]= -1931484818;
assign addr[37190]= -1896833245;
assign addr[37191]= -1859775393;
assign addr[37192]= -1820358275;
assign addr[37193]= -1778631892;
assign addr[37194]= -1734649179;
assign addr[37195]= -1688465931;
assign addr[37196]= -1640140734;
assign addr[37197]= -1589734894;
assign addr[37198]= -1537312353;
assign addr[37199]= -1482939614;
assign addr[37200]= -1426685652;
assign addr[37201]= -1368621831;
assign addr[37202]= -1308821808;
assign addr[37203]= -1247361445;
assign addr[37204]= -1184318708;
assign addr[37205]= -1119773573;
assign addr[37206]= -1053807919;
assign addr[37207]= -986505429;
assign addr[37208]= -917951481;
assign addr[37209]= -848233042;
assign addr[37210]= -777438554;
assign addr[37211]= -705657826;
assign addr[37212]= -632981917;
assign addr[37213]= -559503022;
assign addr[37214]= -485314355;
assign addr[37215]= -410510029;
assign addr[37216]= -335184940;
assign addr[37217]= -259434643;
assign addr[37218]= -183355234;
assign addr[37219]= -107043224;
assign addr[37220]= -30595422;
assign addr[37221]= 45891193;
assign addr[37222]= 122319591;
assign addr[37223]= 198592817;
assign addr[37224]= 274614114;
assign addr[37225]= 350287041;
assign addr[37226]= 425515602;
assign addr[37227]= 500204365;
assign addr[37228]= 574258580;
assign addr[37229]= 647584304;
assign addr[37230]= 720088517;
assign addr[37231]= 791679244;
assign addr[37232]= 862265664;
assign addr[37233]= 931758235;
assign addr[37234]= 1000068799;
assign addr[37235]= 1067110699;
assign addr[37236]= 1132798888;
assign addr[37237]= 1197050035;
assign addr[37238]= 1259782632;
assign addr[37239]= 1320917099;
assign addr[37240]= 1380375881;
assign addr[37241]= 1438083551;
assign addr[37242]= 1493966902;
assign addr[37243]= 1547955041;
assign addr[37244]= 1599979481;
assign addr[37245]= 1649974225;
assign addr[37246]= 1697875851;
assign addr[37247]= 1743623590;
assign addr[37248]= 1787159411;
assign addr[37249]= 1828428082;
assign addr[37250]= 1867377253;
assign addr[37251]= 1903957513;
assign addr[37252]= 1938122457;
assign addr[37253]= 1969828744;
assign addr[37254]= 1999036154;
assign addr[37255]= 2025707632;
assign addr[37256]= 2049809346;
assign addr[37257]= 2071310720;
assign addr[37258]= 2090184478;
assign addr[37259]= 2106406677;
assign addr[37260]= 2119956737;
assign addr[37261]= 2130817471;
assign addr[37262]= 2138975100;
assign addr[37263]= 2144419275;
assign addr[37264]= 2147143090;
assign addr[37265]= 2147143090;
assign addr[37266]= 2144419275;
assign addr[37267]= 2138975100;
assign addr[37268]= 2130817471;
assign addr[37269]= 2119956737;
assign addr[37270]= 2106406677;
assign addr[37271]= 2090184478;
assign addr[37272]= 2071310720;
assign addr[37273]= 2049809346;
assign addr[37274]= 2025707632;
assign addr[37275]= 1999036154;
assign addr[37276]= 1969828744;
assign addr[37277]= 1938122457;
assign addr[37278]= 1903957513;
assign addr[37279]= 1867377253;
assign addr[37280]= 1828428082;
assign addr[37281]= 1787159411;
assign addr[37282]= 1743623590;
assign addr[37283]= 1697875851;
assign addr[37284]= 1649974225;
assign addr[37285]= 1599979481;
assign addr[37286]= 1547955041;
assign addr[37287]= 1493966902;
assign addr[37288]= 1438083551;
assign addr[37289]= 1380375881;
assign addr[37290]= 1320917099;
assign addr[37291]= 1259782632;
assign addr[37292]= 1197050035;
assign addr[37293]= 1132798888;
assign addr[37294]= 1067110699;
assign addr[37295]= 1000068799;
assign addr[37296]= 931758235;
assign addr[37297]= 862265664;
assign addr[37298]= 791679244;
assign addr[37299]= 720088517;
assign addr[37300]= 647584304;
assign addr[37301]= 574258580;
assign addr[37302]= 500204365;
assign addr[37303]= 425515602;
assign addr[37304]= 350287041;
assign addr[37305]= 274614114;
assign addr[37306]= 198592817;
assign addr[37307]= 122319591;
assign addr[37308]= 45891193;
assign addr[37309]= -30595422;
assign addr[37310]= -107043224;
assign addr[37311]= -183355234;
assign addr[37312]= -259434643;
assign addr[37313]= -335184940;
assign addr[37314]= -410510029;
assign addr[37315]= -485314355;
assign addr[37316]= -559503022;
assign addr[37317]= -632981917;
assign addr[37318]= -705657826;
assign addr[37319]= -777438554;
assign addr[37320]= -848233042;
assign addr[37321]= -917951481;
assign addr[37322]= -986505429;
assign addr[37323]= -1053807919;
assign addr[37324]= -1119773573;
assign addr[37325]= -1184318708;
assign addr[37326]= -1247361445;
assign addr[37327]= -1308821808;
assign addr[37328]= -1368621831;
assign addr[37329]= -1426685652;
assign addr[37330]= -1482939614;
assign addr[37331]= -1537312353;
assign addr[37332]= -1589734894;
assign addr[37333]= -1640140734;
assign addr[37334]= -1688465931;
assign addr[37335]= -1734649179;
assign addr[37336]= -1778631892;
assign addr[37337]= -1820358275;
assign addr[37338]= -1859775393;
assign addr[37339]= -1896833245;
assign addr[37340]= -1931484818;
assign addr[37341]= -1963686155;
assign addr[37342]= -1993396407;
assign addr[37343]= -2020577882;
assign addr[37344]= -2045196100;
assign addr[37345]= -2067219829;
assign addr[37346]= -2086621133;
assign addr[37347]= -2103375398;
assign addr[37348]= -2117461370;
assign addr[37349]= -2128861181;
assign addr[37350]= -2137560369;
assign addr[37351]= -2143547897;
assign addr[37352]= -2146816171;
assign addr[37353]= -2147361045;
assign addr[37354]= -2145181827;
assign addr[37355]= -2140281282;
assign addr[37356]= -2132665626;
assign addr[37357]= -2122344521;
assign addr[37358]= -2109331059;
assign addr[37359]= -2093641749;
assign addr[37360]= -2075296495;
assign addr[37361]= -2054318569;
assign addr[37362]= -2030734582;
assign addr[37363]= -2004574453;
assign addr[37364]= -1975871368;
assign addr[37365]= -1944661739;
assign addr[37366]= -1910985158;
assign addr[37367]= -1874884346;
assign addr[37368]= -1836405100;
assign addr[37369]= -1795596234;
assign addr[37370]= -1752509516;
assign addr[37371]= -1707199606;
assign addr[37372]= -1659723983;
assign addr[37373]= -1610142873;
assign addr[37374]= -1558519173;
assign addr[37375]= -1504918373;
assign addr[37376]= -1449408469;
assign addr[37377]= -1392059879;
assign addr[37378]= -1332945355;
assign addr[37379]= -1272139887;
assign addr[37380]= -1209720613;
assign addr[37381]= -1145766716;
assign addr[37382]= -1080359326;
assign addr[37383]= -1013581418;
assign addr[37384]= -945517704;
assign addr[37385]= -876254528;
assign addr[37386]= -805879757;
assign addr[37387]= -734482665;
assign addr[37388]= -662153826;
assign addr[37389]= -588984994;
assign addr[37390]= -515068990;
assign addr[37391]= -440499581;
assign addr[37392]= -365371365;
assign addr[37393]= -289779648;
assign addr[37394]= -213820322;
assign addr[37395]= -137589750;
assign addr[37396]= -61184634;
assign addr[37397]= 15298099;
assign addr[37398]= 91761426;
assign addr[37399]= 168108346;
assign addr[37400]= 244242007;
assign addr[37401]= 320065829;
assign addr[37402]= 395483624;
assign addr[37403]= 470399716;
assign addr[37404]= 544719071;
assign addr[37405]= 618347408;
assign addr[37406]= 691191324;
assign addr[37407]= 763158411;
assign addr[37408]= 834157373;
assign addr[37409]= 904098143;
assign addr[37410]= 972891995;
assign addr[37411]= 1040451659;
assign addr[37412]= 1106691431;
assign addr[37413]= 1171527280;
assign addr[37414]= 1234876957;
assign addr[37415]= 1296660098;
assign addr[37416]= 1356798326;
assign addr[37417]= 1415215352;
assign addr[37418]= 1471837070;
assign addr[37419]= 1526591649;
assign addr[37420]= 1579409630;
assign addr[37421]= 1630224009;
assign addr[37422]= 1678970324;
assign addr[37423]= 1725586737;
assign addr[37424]= 1770014111;
assign addr[37425]= 1812196087;
assign addr[37426]= 1852079154;
assign addr[37427]= 1889612716;
assign addr[37428]= 1924749160;
assign addr[37429]= 1957443913;
assign addr[37430]= 1987655498;
assign addr[37431]= 2015345591;
assign addr[37432]= 2040479063;
assign addr[37433]= 2063024031;
assign addr[37434]= 2082951896;
assign addr[37435]= 2100237377;
assign addr[37436]= 2114858546;
assign addr[37437]= 2126796855;
assign addr[37438]= 2136037160;
assign addr[37439]= 2142567738;
assign addr[37440]= 2146380306;
assign addr[37441]= 2147470025;
assign addr[37442]= 2145835515;
assign addr[37443]= 2141478848;
assign addr[37444]= 2134405552;
assign addr[37445]= 2124624598;
assign addr[37446]= 2112148396;
assign addr[37447]= 2096992772;
assign addr[37448]= 2079176953;
assign addr[37449]= 2058723538;
assign addr[37450]= 2035658475;
assign addr[37451]= 2010011024;
assign addr[37452]= 1981813720;
assign addr[37453]= 1951102334;
assign addr[37454]= 1917915825;
assign addr[37455]= 1882296293;
assign addr[37456]= 1844288924;
assign addr[37457]= 1803941934;
assign addr[37458]= 1761306505;
assign addr[37459]= 1716436725;
assign addr[37460]= 1669389513;
assign addr[37461]= 1620224553;
assign addr[37462]= 1569004214;
assign addr[37463]= 1515793473;
assign addr[37464]= 1460659832;
assign addr[37465]= 1403673233;
assign addr[37466]= 1344905966;
assign addr[37467]= 1284432584;
assign addr[37468]= 1222329801;
assign addr[37469]= 1158676398;
assign addr[37470]= 1093553126;
assign addr[37471]= 1027042599;
assign addr[37472]= 959229189;
assign addr[37473]= 890198924;
assign addr[37474]= 820039373;
assign addr[37475]= 748839539;
assign addr[37476]= 676689746;
assign addr[37477]= 603681519;
assign addr[37478]= 529907477;
assign addr[37479]= 455461206;
assign addr[37480]= 380437148;
assign addr[37481]= 304930476;
assign addr[37482]= 229036977;
assign addr[37483]= 152852926;
assign addr[37484]= 76474970;
assign addr[37485]= 0;
assign addr[37486]= -76474970;
assign addr[37487]= -152852926;
assign addr[37488]= -229036977;
assign addr[37489]= -304930476;
assign addr[37490]= -380437148;
assign addr[37491]= -455461206;
assign addr[37492]= -529907477;
assign addr[37493]= -603681519;
assign addr[37494]= -676689746;
assign addr[37495]= -748839539;
assign addr[37496]= -820039373;
assign addr[37497]= -890198924;
assign addr[37498]= -959229189;
assign addr[37499]= -1027042599;
assign addr[37500]= -1093553126;
assign addr[37501]= -1158676398;
assign addr[37502]= -1222329801;
assign addr[37503]= -1284432584;
assign addr[37504]= -1344905966;
assign addr[37505]= -1403673233;
assign addr[37506]= -1460659832;
assign addr[37507]= -1515793473;
assign addr[37508]= -1569004214;
assign addr[37509]= -1620224553;
assign addr[37510]= -1669389513;
assign addr[37511]= -1716436725;
assign addr[37512]= -1761306505;
assign addr[37513]= -1803941934;
assign addr[37514]= -1844288924;
assign addr[37515]= -1882296293;
assign addr[37516]= -1917915825;
assign addr[37517]= -1951102334;
assign addr[37518]= -1981813720;
assign addr[37519]= -2010011024;
assign addr[37520]= -2035658475;
assign addr[37521]= -2058723538;
assign addr[37522]= -2079176953;
assign addr[37523]= -2096992772;
assign addr[37524]= -2112148396;
assign addr[37525]= -2124624598;
assign addr[37526]= -2134405552;
assign addr[37527]= -2141478848;
assign addr[37528]= -2145835515;
assign addr[37529]= -2147470025;
assign addr[37530]= -2146380306;
assign addr[37531]= -2142567738;
assign addr[37532]= -2136037160;
assign addr[37533]= -2126796855;
assign addr[37534]= -2114858546;
assign addr[37535]= -2100237377;
assign addr[37536]= -2082951896;
assign addr[37537]= -2063024031;
assign addr[37538]= -2040479063;
assign addr[37539]= -2015345591;
assign addr[37540]= -1987655498;
assign addr[37541]= -1957443913;
assign addr[37542]= -1924749160;
assign addr[37543]= -1889612716;
assign addr[37544]= -1852079154;
assign addr[37545]= -1812196087;
assign addr[37546]= -1770014111;
assign addr[37547]= -1725586737;
assign addr[37548]= -1678970324;
assign addr[37549]= -1630224009;
assign addr[37550]= -1579409630;
assign addr[37551]= -1526591649;
assign addr[37552]= -1471837070;
assign addr[37553]= -1415215352;
assign addr[37554]= -1356798326;
assign addr[37555]= -1296660098;
assign addr[37556]= -1234876957;
assign addr[37557]= -1171527280;
assign addr[37558]= -1106691431;
assign addr[37559]= -1040451659;
assign addr[37560]= -972891995;
assign addr[37561]= -904098143;
assign addr[37562]= -834157373;
assign addr[37563]= -763158411;
assign addr[37564]= -691191324;
assign addr[37565]= -618347408;
assign addr[37566]= -544719071;
assign addr[37567]= -470399716;
assign addr[37568]= -395483624;
assign addr[37569]= -320065829;
assign addr[37570]= -244242007;
assign addr[37571]= -168108346;
assign addr[37572]= -91761426;
assign addr[37573]= -15298099;
assign addr[37574]= 61184634;
assign addr[37575]= 137589750;
assign addr[37576]= 213820322;
assign addr[37577]= 289779648;
assign addr[37578]= 365371365;
assign addr[37579]= 440499581;
assign addr[37580]= 515068990;
assign addr[37581]= 588984994;
assign addr[37582]= 662153826;
assign addr[37583]= 734482665;
assign addr[37584]= 805879757;
assign addr[37585]= 876254528;
assign addr[37586]= 945517704;
assign addr[37587]= 1013581418;
assign addr[37588]= 1080359326;
assign addr[37589]= 1145766716;
assign addr[37590]= 1209720613;
assign addr[37591]= 1272139887;
assign addr[37592]= 1332945355;
assign addr[37593]= 1392059879;
assign addr[37594]= 1449408469;
assign addr[37595]= 1504918373;
assign addr[37596]= 1558519173;
assign addr[37597]= 1610142873;
assign addr[37598]= 1659723983;
assign addr[37599]= 1707199606;
assign addr[37600]= 1752509516;
assign addr[37601]= 1795596234;
assign addr[37602]= 1836405100;
assign addr[37603]= 1874884346;
assign addr[37604]= 1910985158;
assign addr[37605]= 1944661739;
assign addr[37606]= 1975871368;
assign addr[37607]= 2004574453;
assign addr[37608]= 2030734582;
assign addr[37609]= 2054318569;
assign addr[37610]= 2075296495;
assign addr[37611]= 2093641749;
assign addr[37612]= 2109331059;
assign addr[37613]= 2122344521;
assign addr[37614]= 2132665626;
assign addr[37615]= 2140281282;
assign addr[37616]= 2145181827;
assign addr[37617]= 2147361045;
assign addr[37618]= 2146816171;
assign addr[37619]= 2143547897;
assign addr[37620]= 2137560369;
assign addr[37621]= 2128861181;
assign addr[37622]= 2117461370;
assign addr[37623]= 2103375398;
assign addr[37624]= 2086621133;
assign addr[37625]= 2067219829;
assign addr[37626]= 2045196100;
assign addr[37627]= 2020577882;
assign addr[37628]= 1993396407;
assign addr[37629]= 1963686155;
assign addr[37630]= 1931484818;
assign addr[37631]= 1896833245;
assign addr[37632]= 1859775393;
assign addr[37633]= 1820358275;
assign addr[37634]= 1778631892;
assign addr[37635]= 1734649179;
assign addr[37636]= 1688465931;
assign addr[37637]= 1640140734;
assign addr[37638]= 1589734894;
assign addr[37639]= 1537312353;
assign addr[37640]= 1482939614;
assign addr[37641]= 1426685652;
assign addr[37642]= 1368621831;
assign addr[37643]= 1308821808;
assign addr[37644]= 1247361445;
assign addr[37645]= 1184318708;
assign addr[37646]= 1119773573;
assign addr[37647]= 1053807919;
assign addr[37648]= 986505429;
assign addr[37649]= 917951481;
assign addr[37650]= 848233042;
assign addr[37651]= 777438554;
assign addr[37652]= 705657826;
assign addr[37653]= 632981917;
assign addr[37654]= 559503022;
assign addr[37655]= 485314355;
assign addr[37656]= 410510029;
assign addr[37657]= 335184940;
assign addr[37658]= 259434643;
assign addr[37659]= 183355234;
assign addr[37660]= 107043224;
assign addr[37661]= 30595422;
assign addr[37662]= -45891193;
assign addr[37663]= -122319591;
assign addr[37664]= -198592817;
assign addr[37665]= -274614114;
assign addr[37666]= -350287041;
assign addr[37667]= -425515602;
assign addr[37668]= -500204365;
assign addr[37669]= -574258580;
assign addr[37670]= -647584304;
assign addr[37671]= -720088517;
assign addr[37672]= -791679244;
assign addr[37673]= -862265664;
assign addr[37674]= -931758235;
assign addr[37675]= -1000068799;
assign addr[37676]= -1067110699;
assign addr[37677]= -1132798888;
assign addr[37678]= -1197050035;
assign addr[37679]= -1259782632;
assign addr[37680]= -1320917099;
assign addr[37681]= -1380375881;
assign addr[37682]= -1438083551;
assign addr[37683]= -1493966902;
assign addr[37684]= -1547955041;
assign addr[37685]= -1599979481;
assign addr[37686]= -1649974225;
assign addr[37687]= -1697875851;
assign addr[37688]= -1743623590;
assign addr[37689]= -1787159411;
assign addr[37690]= -1828428082;
assign addr[37691]= -1867377253;
assign addr[37692]= -1903957513;
assign addr[37693]= -1938122457;
assign addr[37694]= -1969828744;
assign addr[37695]= -1999036154;
assign addr[37696]= -2025707632;
assign addr[37697]= -2049809346;
assign addr[37698]= -2071310720;
assign addr[37699]= -2090184478;
assign addr[37700]= -2106406677;
assign addr[37701]= -2119956737;
assign addr[37702]= -2130817471;
assign addr[37703]= -2138975100;
assign addr[37704]= -2144419275;
assign addr[37705]= -2147143090;
assign addr[37706]= -2147143090;
assign addr[37707]= -2144419275;
assign addr[37708]= -2138975100;
assign addr[37709]= -2130817471;
assign addr[37710]= -2119956737;
assign addr[37711]= -2106406677;
assign addr[37712]= -2090184478;
assign addr[37713]= -2071310720;
assign addr[37714]= -2049809346;
assign addr[37715]= -2025707632;
assign addr[37716]= -1999036154;
assign addr[37717]= -1969828744;
assign addr[37718]= -1938122457;
assign addr[37719]= -1903957513;
assign addr[37720]= -1867377253;
assign addr[37721]= -1828428082;
assign addr[37722]= -1787159411;
assign addr[37723]= -1743623590;
assign addr[37724]= -1697875851;
assign addr[37725]= -1649974225;
assign addr[37726]= -1599979481;
assign addr[37727]= -1547955041;
assign addr[37728]= -1493966902;
assign addr[37729]= -1438083551;
assign addr[37730]= -1380375881;
assign addr[37731]= -1320917099;
assign addr[37732]= -1259782632;
assign addr[37733]= -1197050035;
assign addr[37734]= -1132798888;
assign addr[37735]= -1067110699;
assign addr[37736]= -1000068799;
assign addr[37737]= -931758235;
assign addr[37738]= -862265664;
assign addr[37739]= -791679244;
assign addr[37740]= -720088517;
assign addr[37741]= -647584304;
assign addr[37742]= -574258580;
assign addr[37743]= -500204365;
assign addr[37744]= -425515602;
assign addr[37745]= -350287041;
assign addr[37746]= -274614114;
assign addr[37747]= -198592817;
assign addr[37748]= -122319591;
assign addr[37749]= -45891193;
assign addr[37750]= 30595422;
assign addr[37751]= 107043224;
assign addr[37752]= 183355234;
assign addr[37753]= 259434643;
assign addr[37754]= 335184940;
assign addr[37755]= 410510029;
assign addr[37756]= 485314355;
assign addr[37757]= 559503022;
assign addr[37758]= 632981917;
assign addr[37759]= 705657826;
assign addr[37760]= 777438554;
assign addr[37761]= 848233042;
assign addr[37762]= 917951481;
assign addr[37763]= 986505429;
assign addr[37764]= 1053807919;
assign addr[37765]= 1119773573;
assign addr[37766]= 1184318708;
assign addr[37767]= 1247361445;
assign addr[37768]= 1308821808;
assign addr[37769]= 1368621831;
assign addr[37770]= 1426685652;
assign addr[37771]= 1482939614;
assign addr[37772]= 1537312353;
assign addr[37773]= 1589734894;
assign addr[37774]= 1640140734;
assign addr[37775]= 1688465931;
assign addr[37776]= 1734649179;
assign addr[37777]= 1778631892;
assign addr[37778]= 1820358275;
assign addr[37779]= 1859775393;
assign addr[37780]= 1896833245;
assign addr[37781]= 1931484818;
assign addr[37782]= 1963686155;
assign addr[37783]= 1993396407;
assign addr[37784]= 2020577882;
assign addr[37785]= 2045196100;
assign addr[37786]= 2067219829;
assign addr[37787]= 2086621133;
assign addr[37788]= 2103375398;
assign addr[37789]= 2117461370;
assign addr[37790]= 2128861181;
assign addr[37791]= 2137560369;
assign addr[37792]= 2143547897;
assign addr[37793]= 2146816171;
assign addr[37794]= 2147361045;
assign addr[37795]= 2145181827;
assign addr[37796]= 2140281282;
assign addr[37797]= 2132665626;
assign addr[37798]= 2122344521;
assign addr[37799]= 2109331059;
assign addr[37800]= 2093641749;
assign addr[37801]= 2075296495;
assign addr[37802]= 2054318569;
assign addr[37803]= 2030734582;
assign addr[37804]= 2004574453;
assign addr[37805]= 1975871368;
assign addr[37806]= 1944661739;
assign addr[37807]= 1910985158;
assign addr[37808]= 1874884346;
assign addr[37809]= 1836405100;
assign addr[37810]= 1795596234;
assign addr[37811]= 1752509516;
assign addr[37812]= 1707199606;
assign addr[37813]= 1659723983;
assign addr[37814]= 1610142873;
assign addr[37815]= 1558519173;
assign addr[37816]= 1504918373;
assign addr[37817]= 1449408469;
assign addr[37818]= 1392059879;
assign addr[37819]= 1332945355;
assign addr[37820]= 1272139887;
assign addr[37821]= 1209720613;
assign addr[37822]= 1145766716;
assign addr[37823]= 1080359326;
assign addr[37824]= 1013581418;
assign addr[37825]= 945517704;
assign addr[37826]= 876254528;
assign addr[37827]= 805879757;
assign addr[37828]= 734482665;
assign addr[37829]= 662153826;
assign addr[37830]= 588984994;
assign addr[37831]= 515068990;
assign addr[37832]= 440499581;
assign addr[37833]= 365371365;
assign addr[37834]= 289779648;
assign addr[37835]= 213820322;
assign addr[37836]= 137589750;
assign addr[37837]= 61184634;
assign addr[37838]= -15298099;
assign addr[37839]= -91761426;
assign addr[37840]= -168108346;
assign addr[37841]= -244242007;
assign addr[37842]= -320065829;
assign addr[37843]= -395483624;
assign addr[37844]= -470399716;
assign addr[37845]= -544719071;
assign addr[37846]= -618347408;
assign addr[37847]= -691191324;
assign addr[37848]= -763158411;
assign addr[37849]= -834157373;
assign addr[37850]= -904098143;
assign addr[37851]= -972891995;
assign addr[37852]= -1040451659;
assign addr[37853]= -1106691431;
assign addr[37854]= -1171527280;
assign addr[37855]= -1234876957;
assign addr[37856]= -1296660098;
assign addr[37857]= -1356798326;
assign addr[37858]= -1415215352;
assign addr[37859]= -1471837070;
assign addr[37860]= -1526591649;
assign addr[37861]= -1579409630;
assign addr[37862]= -1630224009;
assign addr[37863]= -1678970324;
assign addr[37864]= -1725586737;
assign addr[37865]= -1770014111;
assign addr[37866]= -1812196087;
assign addr[37867]= -1852079154;
assign addr[37868]= -1889612716;
assign addr[37869]= -1924749160;
assign addr[37870]= -1957443913;
assign addr[37871]= -1987655498;
assign addr[37872]= -2015345591;
assign addr[37873]= -2040479063;
assign addr[37874]= -2063024031;
assign addr[37875]= -2082951896;
assign addr[37876]= -2100237377;
assign addr[37877]= -2114858546;
assign addr[37878]= -2126796855;
assign addr[37879]= -2136037160;
assign addr[37880]= -2142567738;
assign addr[37881]= -2146380306;
assign addr[37882]= -2147470025;
assign addr[37883]= -2145835515;
assign addr[37884]= -2141478848;
assign addr[37885]= -2134405552;
assign addr[37886]= -2124624598;
assign addr[37887]= -2112148396;
assign addr[37888]= -2096992772;
assign addr[37889]= -2079176953;
assign addr[37890]= -2058723538;
assign addr[37891]= -2035658475;
assign addr[37892]= -2010011024;
assign addr[37893]= -1981813720;
assign addr[37894]= -1951102334;
assign addr[37895]= -1917915825;
assign addr[37896]= -1882296293;
assign addr[37897]= -1844288924;
assign addr[37898]= -1803941934;
assign addr[37899]= -1761306505;
assign addr[37900]= -1716436725;
assign addr[37901]= -1669389513;
assign addr[37902]= -1620224553;
assign addr[37903]= -1569004214;
assign addr[37904]= -1515793473;
assign addr[37905]= -1460659832;
assign addr[37906]= -1403673233;
assign addr[37907]= -1344905966;
assign addr[37908]= -1284432584;
assign addr[37909]= -1222329801;
assign addr[37910]= -1158676398;
assign addr[37911]= -1093553126;
assign addr[37912]= -1027042599;
assign addr[37913]= -959229189;
assign addr[37914]= -890198924;
assign addr[37915]= -820039373;
assign addr[37916]= -748839539;
assign addr[37917]= -676689746;
assign addr[37918]= -603681519;
assign addr[37919]= -529907477;
assign addr[37920]= -455461206;
assign addr[37921]= -380437148;
assign addr[37922]= -304930476;
assign addr[37923]= -229036977;
assign addr[37924]= -152852926;
assign addr[37925]= -76474970;
assign addr[37926]= 0;
assign addr[37927]= 76474970;
assign addr[37928]= 152852926;
assign addr[37929]= 229036977;
assign addr[37930]= 304930476;
assign addr[37931]= 380437148;
assign addr[37932]= 455461206;
assign addr[37933]= 529907477;
assign addr[37934]= 603681519;
assign addr[37935]= 676689746;
assign addr[37936]= 748839539;
assign addr[37937]= 820039373;
assign addr[37938]= 890198924;
assign addr[37939]= 959229189;
assign addr[37940]= 1027042599;
assign addr[37941]= 1093553126;
assign addr[37942]= 1158676398;
assign addr[37943]= 1222329801;
assign addr[37944]= 1284432584;
assign addr[37945]= 1344905966;
assign addr[37946]= 1403673233;
assign addr[37947]= 1460659832;
assign addr[37948]= 1515793473;
assign addr[37949]= 1569004214;
assign addr[37950]= 1620224553;
assign addr[37951]= 1669389513;
assign addr[37952]= 1716436725;
assign addr[37953]= 1761306505;
assign addr[37954]= 1803941934;
assign addr[37955]= 1844288924;
assign addr[37956]= 1882296293;
assign addr[37957]= 1917915825;
assign addr[37958]= 1951102334;
assign addr[37959]= 1981813720;
assign addr[37960]= 2010011024;
assign addr[37961]= 2035658475;
assign addr[37962]= 2058723538;
assign addr[37963]= 2079176953;
assign addr[37964]= 2096992772;
assign addr[37965]= 2112148396;
assign addr[37966]= 2124624598;
assign addr[37967]= 2134405552;
assign addr[37968]= 2141478848;
assign addr[37969]= 2145835515;
assign addr[37970]= 2147470025;
assign addr[37971]= 2146380306;
assign addr[37972]= 2142567738;
assign addr[37973]= 2136037160;
assign addr[37974]= 2126796855;
assign addr[37975]= 2114858546;
assign addr[37976]= 2100237377;
assign addr[37977]= 2082951896;
assign addr[37978]= 2063024031;
assign addr[37979]= 2040479063;
assign addr[37980]= 2015345591;
assign addr[37981]= 1987655498;
assign addr[37982]= 1957443913;
assign addr[37983]= 1924749160;
assign addr[37984]= 1889612716;
assign addr[37985]= 1852079154;
assign addr[37986]= 1812196087;
assign addr[37987]= 1770014111;
assign addr[37988]= 1725586737;
assign addr[37989]= 1678970324;
assign addr[37990]= 1630224009;
assign addr[37991]= 1579409630;
assign addr[37992]= 1526591649;
assign addr[37993]= 1471837070;
assign addr[37994]= 1415215352;
assign addr[37995]= 1356798326;
assign addr[37996]= 1296660098;
assign addr[37997]= 1234876957;
assign addr[37998]= 1171527280;
assign addr[37999]= 1106691431;
assign addr[38000]= 1040451659;
assign addr[38001]= 972891995;
assign addr[38002]= 904098143;
assign addr[38003]= 834157373;
assign addr[38004]= 763158411;
assign addr[38005]= 691191324;
assign addr[38006]= 618347408;
assign addr[38007]= 544719071;
assign addr[38008]= 470399716;
assign addr[38009]= 395483624;
assign addr[38010]= 320065829;
assign addr[38011]= 244242007;
assign addr[38012]= 168108346;
assign addr[38013]= 91761426;
assign addr[38014]= 15298099;
assign addr[38015]= -61184634;
assign addr[38016]= -137589750;
assign addr[38017]= -213820322;
assign addr[38018]= -289779648;
assign addr[38019]= -365371365;
assign addr[38020]= -440499581;
assign addr[38021]= -515068990;
assign addr[38022]= -588984994;
assign addr[38023]= -662153826;
assign addr[38024]= -734482665;
assign addr[38025]= -805879757;
assign addr[38026]= -876254528;
assign addr[38027]= -945517704;
assign addr[38028]= -1013581418;
assign addr[38029]= -1080359326;
assign addr[38030]= -1145766716;
assign addr[38031]= -1209720613;
assign addr[38032]= -1272139887;
assign addr[38033]= -1332945355;
assign addr[38034]= -1392059879;
assign addr[38035]= -1449408469;
assign addr[38036]= -1504918373;
assign addr[38037]= -1558519173;
assign addr[38038]= -1610142873;
assign addr[38039]= -1659723983;
assign addr[38040]= -1707199606;
assign addr[38041]= -1752509516;
assign addr[38042]= -1795596234;
assign addr[38043]= -1836405100;
assign addr[38044]= -1874884346;
assign addr[38045]= -1910985158;
assign addr[38046]= -1944661739;
assign addr[38047]= -1975871368;
assign addr[38048]= -2004574453;
assign addr[38049]= -2030734582;
assign addr[38050]= -2054318569;
assign addr[38051]= -2075296495;
assign addr[38052]= -2093641749;
assign addr[38053]= -2109331059;
assign addr[38054]= -2122344521;
assign addr[38055]= -2132665626;
assign addr[38056]= -2140281282;
assign addr[38057]= -2145181827;
assign addr[38058]= -2147361045;
assign addr[38059]= -2146816171;
assign addr[38060]= -2143547897;
assign addr[38061]= -2137560369;
assign addr[38062]= -2128861181;
assign addr[38063]= -2117461370;
assign addr[38064]= -2103375398;
assign addr[38065]= -2086621133;
assign addr[38066]= -2067219829;
assign addr[38067]= -2045196100;
assign addr[38068]= -2020577882;
assign addr[38069]= -1993396407;
assign addr[38070]= -1963686155;
assign addr[38071]= -1931484818;
assign addr[38072]= -1896833245;
assign addr[38073]= -1859775393;
assign addr[38074]= -1820358275;
assign addr[38075]= -1778631892;
assign addr[38076]= -1734649179;
assign addr[38077]= -1688465931;
assign addr[38078]= -1640140734;
assign addr[38079]= -1589734894;
assign addr[38080]= -1537312353;
assign addr[38081]= -1482939614;
assign addr[38082]= -1426685652;
assign addr[38083]= -1368621831;
assign addr[38084]= -1308821808;
assign addr[38085]= -1247361445;
assign addr[38086]= -1184318708;
assign addr[38087]= -1119773573;
assign addr[38088]= -1053807919;
assign addr[38089]= -986505429;
assign addr[38090]= -917951481;
assign addr[38091]= -848233042;
assign addr[38092]= -777438554;
assign addr[38093]= -705657826;
assign addr[38094]= -632981917;
assign addr[38095]= -559503022;
assign addr[38096]= -485314355;
assign addr[38097]= -410510029;
assign addr[38098]= -335184940;
assign addr[38099]= -259434643;
assign addr[38100]= -183355234;
assign addr[38101]= -107043224;
assign addr[38102]= -30595422;
assign addr[38103]= 45891193;
assign addr[38104]= 122319591;
assign addr[38105]= 198592817;
assign addr[38106]= 274614114;
assign addr[38107]= 350287041;
assign addr[38108]= 425515602;
assign addr[38109]= 500204365;
assign addr[38110]= 574258580;
assign addr[38111]= 647584304;
assign addr[38112]= 720088517;
assign addr[38113]= 791679244;
assign addr[38114]= 862265664;
assign addr[38115]= 931758235;
assign addr[38116]= 1000068799;
assign addr[38117]= 1067110699;
assign addr[38118]= 1132798888;
assign addr[38119]= 1197050035;
assign addr[38120]= 1259782632;
assign addr[38121]= 1320917099;
assign addr[38122]= 1380375881;
assign addr[38123]= 1438083551;
assign addr[38124]= 1493966902;
assign addr[38125]= 1547955041;
assign addr[38126]= 1599979481;
assign addr[38127]= 1649974225;
assign addr[38128]= 1697875851;
assign addr[38129]= 1743623590;
assign addr[38130]= 1787159411;
assign addr[38131]= 1828428082;
assign addr[38132]= 1867377253;
assign addr[38133]= 1903957513;
assign addr[38134]= 1938122457;
assign addr[38135]= 1969828744;
assign addr[38136]= 1999036154;
assign addr[38137]= 2025707632;
assign addr[38138]= 2049809346;
assign addr[38139]= 2071310720;
assign addr[38140]= 2090184478;
assign addr[38141]= 2106406677;
assign addr[38142]= 2119956737;
assign addr[38143]= 2130817471;
assign addr[38144]= 2138975100;
assign addr[38145]= 2144419275;
assign addr[38146]= 2147143090;
assign addr[38147]= 2147143090;
assign addr[38148]= 2144419275;
assign addr[38149]= 2138975100;
assign addr[38150]= 2130817471;
assign addr[38151]= 2119956737;
assign addr[38152]= 2106406677;
assign addr[38153]= 2090184478;
assign addr[38154]= 2071310720;
assign addr[38155]= 2049809346;
assign addr[38156]= 2025707632;
assign addr[38157]= 1999036154;
assign addr[38158]= 1969828744;
assign addr[38159]= 1938122457;
assign addr[38160]= 1903957513;
assign addr[38161]= 1867377253;
assign addr[38162]= 1828428082;
assign addr[38163]= 1787159411;
assign addr[38164]= 1743623590;
assign addr[38165]= 1697875851;
assign addr[38166]= 1649974225;
assign addr[38167]= 1599979481;
assign addr[38168]= 1547955041;
assign addr[38169]= 1493966902;
assign addr[38170]= 1438083551;
assign addr[38171]= 1380375881;
assign addr[38172]= 1320917099;
assign addr[38173]= 1259782632;
assign addr[38174]= 1197050035;
assign addr[38175]= 1132798888;
assign addr[38176]= 1067110699;
assign addr[38177]= 1000068799;
assign addr[38178]= 931758235;
assign addr[38179]= 862265664;
assign addr[38180]= 791679244;
assign addr[38181]= 720088517;
assign addr[38182]= 647584304;
assign addr[38183]= 574258580;
assign addr[38184]= 500204365;
assign addr[38185]= 425515602;
assign addr[38186]= 350287041;
assign addr[38187]= 274614114;
assign addr[38188]= 198592817;
assign addr[38189]= 122319591;
assign addr[38190]= 45891193;
assign addr[38191]= -30595422;
assign addr[38192]= -107043224;
assign addr[38193]= -183355234;
assign addr[38194]= -259434643;
assign addr[38195]= -335184940;
assign addr[38196]= -410510029;
assign addr[38197]= -485314355;
assign addr[38198]= -559503022;
assign addr[38199]= -632981917;
assign addr[38200]= -705657826;
assign addr[38201]= -777438554;
assign addr[38202]= -848233042;
assign addr[38203]= -917951481;
assign addr[38204]= -986505429;
assign addr[38205]= -1053807919;
assign addr[38206]= -1119773573;
assign addr[38207]= -1184318708;
assign addr[38208]= -1247361445;
assign addr[38209]= -1308821808;
assign addr[38210]= -1368621831;
assign addr[38211]= -1426685652;
assign addr[38212]= -1482939614;
assign addr[38213]= -1537312353;
assign addr[38214]= -1589734894;
assign addr[38215]= -1640140734;
assign addr[38216]= -1688465931;
assign addr[38217]= -1734649179;
assign addr[38218]= -1778631892;
assign addr[38219]= -1820358275;
assign addr[38220]= -1859775393;
assign addr[38221]= -1896833245;
assign addr[38222]= -1931484818;
assign addr[38223]= -1963686155;
assign addr[38224]= -1993396407;
assign addr[38225]= -2020577882;
assign addr[38226]= -2045196100;
assign addr[38227]= -2067219829;
assign addr[38228]= -2086621133;
assign addr[38229]= -2103375398;
assign addr[38230]= -2117461370;
assign addr[38231]= -2128861181;
assign addr[38232]= -2137560369;
assign addr[38233]= -2143547897;
assign addr[38234]= -2146816171;
assign addr[38235]= -2147361045;
assign addr[38236]= -2145181827;
assign addr[38237]= -2140281282;
assign addr[38238]= -2132665626;
assign addr[38239]= -2122344521;
assign addr[38240]= -2109331059;
assign addr[38241]= -2093641749;
assign addr[38242]= -2075296495;
assign addr[38243]= -2054318569;
assign addr[38244]= -2030734582;
assign addr[38245]= -2004574453;
assign addr[38246]= -1975871368;
assign addr[38247]= -1944661739;
assign addr[38248]= -1910985158;
assign addr[38249]= -1874884346;
assign addr[38250]= -1836405100;
assign addr[38251]= -1795596234;
assign addr[38252]= -1752509516;
assign addr[38253]= -1707199606;
assign addr[38254]= -1659723983;
assign addr[38255]= -1610142873;
assign addr[38256]= -1558519173;
assign addr[38257]= -1504918373;
assign addr[38258]= -1449408469;
assign addr[38259]= -1392059879;
assign addr[38260]= -1332945355;
assign addr[38261]= -1272139887;
assign addr[38262]= -1209720613;
assign addr[38263]= -1145766716;
assign addr[38264]= -1080359326;
assign addr[38265]= -1013581418;
assign addr[38266]= -945517704;
assign addr[38267]= -876254528;
assign addr[38268]= -805879757;
assign addr[38269]= -734482665;
assign addr[38270]= -662153826;
assign addr[38271]= -588984994;
assign addr[38272]= -515068990;
assign addr[38273]= -440499581;
assign addr[38274]= -365371365;
assign addr[38275]= -289779648;
assign addr[38276]= -213820322;
assign addr[38277]= -137589750;
assign addr[38278]= -61184634;
assign addr[38279]= 15298099;
assign addr[38280]= 91761426;
assign addr[38281]= 168108346;
assign addr[38282]= 244242007;
assign addr[38283]= 320065829;
assign addr[38284]= 395483624;
assign addr[38285]= 470399716;
assign addr[38286]= 544719071;
assign addr[38287]= 618347408;
assign addr[38288]= 691191324;
assign addr[38289]= 763158411;
assign addr[38290]= 834157373;
assign addr[38291]= 904098143;
assign addr[38292]= 972891995;
assign addr[38293]= 1040451659;
assign addr[38294]= 1106691431;
assign addr[38295]= 1171527280;
assign addr[38296]= 1234876957;
assign addr[38297]= 1296660098;
assign addr[38298]= 1356798326;
assign addr[38299]= 1415215352;
assign addr[38300]= 1471837070;
assign addr[38301]= 1526591649;
assign addr[38302]= 1579409630;
assign addr[38303]= 1630224009;
assign addr[38304]= 1678970324;
assign addr[38305]= 1725586737;
assign addr[38306]= 1770014111;
assign addr[38307]= 1812196087;
assign addr[38308]= 1852079154;
assign addr[38309]= 1889612716;
assign addr[38310]= 1924749160;
assign addr[38311]= 1957443913;
assign addr[38312]= 1987655498;
assign addr[38313]= 2015345591;
assign addr[38314]= 2040479063;
assign addr[38315]= 2063024031;
assign addr[38316]= 2082951896;
assign addr[38317]= 2100237377;
assign addr[38318]= 2114858546;
assign addr[38319]= 2126796855;
assign addr[38320]= 2136037160;
assign addr[38321]= 2142567738;
assign addr[38322]= 2146380306;
assign addr[38323]= 2147470025;
assign addr[38324]= 2145835515;
assign addr[38325]= 2141478848;
assign addr[38326]= 2134405552;
assign addr[38327]= 2124624598;
assign addr[38328]= 2112148396;
assign addr[38329]= 2096992772;
assign addr[38330]= 2079176953;
assign addr[38331]= 2058723538;
assign addr[38332]= 2035658475;
assign addr[38333]= 2010011024;
assign addr[38334]= 1981813720;
assign addr[38335]= 1951102334;
assign addr[38336]= 1917915825;
assign addr[38337]= 1882296293;
assign addr[38338]= 1844288924;
assign addr[38339]= 1803941934;
assign addr[38340]= 1761306505;
assign addr[38341]= 1716436725;
assign addr[38342]= 1669389513;
assign addr[38343]= 1620224553;
assign addr[38344]= 1569004214;
assign addr[38345]= 1515793473;
assign addr[38346]= 1460659832;
assign addr[38347]= 1403673233;
assign addr[38348]= 1344905966;
assign addr[38349]= 1284432584;
assign addr[38350]= 1222329801;
assign addr[38351]= 1158676398;
assign addr[38352]= 1093553126;
assign addr[38353]= 1027042599;
assign addr[38354]= 959229189;
assign addr[38355]= 890198924;
assign addr[38356]= 820039373;
assign addr[38357]= 748839539;
assign addr[38358]= 676689746;
assign addr[38359]= 603681519;
assign addr[38360]= 529907477;
assign addr[38361]= 455461206;
assign addr[38362]= 380437148;
assign addr[38363]= 304930476;
assign addr[38364]= 229036977;
assign addr[38365]= 152852926;
assign addr[38366]= 76474970;
assign addr[38367]= 0;
assign addr[38368]= -76474970;
assign addr[38369]= -152852926;
assign addr[38370]= -229036977;
assign addr[38371]= -304930476;
assign addr[38372]= -380437148;
assign addr[38373]= -455461206;
assign addr[38374]= -529907477;
assign addr[38375]= -603681519;
assign addr[38376]= -676689746;
assign addr[38377]= -748839539;
assign addr[38378]= -820039373;
assign addr[38379]= -890198924;
assign addr[38380]= -959229189;
assign addr[38381]= -1027042599;
assign addr[38382]= -1093553126;
assign addr[38383]= -1158676398;
assign addr[38384]= -1222329801;
assign addr[38385]= -1284432584;
assign addr[38386]= -1344905966;
assign addr[38387]= -1403673233;
assign addr[38388]= -1460659832;
assign addr[38389]= -1515793473;
assign addr[38390]= -1569004214;
assign addr[38391]= -1620224553;
assign addr[38392]= -1669389513;
assign addr[38393]= -1716436725;
assign addr[38394]= -1761306505;
assign addr[38395]= -1803941934;
assign addr[38396]= -1844288924;
assign addr[38397]= -1882296293;
assign addr[38398]= -1917915825;
assign addr[38399]= -1951102334;
assign addr[38400]= -1981813720;
assign addr[38401]= -2010011024;
assign addr[38402]= -2035658475;
assign addr[38403]= -2058723538;
assign addr[38404]= -2079176953;
assign addr[38405]= -2096992772;
assign addr[38406]= -2112148396;
assign addr[38407]= -2124624598;
assign addr[38408]= -2134405552;
assign addr[38409]= -2141478848;
assign addr[38410]= -2145835515;
assign addr[38411]= -2147470025;
assign addr[38412]= -2146380306;
assign addr[38413]= -2142567738;
assign addr[38414]= -2136037160;
assign addr[38415]= -2126796855;
assign addr[38416]= -2114858546;
assign addr[38417]= -2100237377;
assign addr[38418]= -2082951896;
assign addr[38419]= -2063024031;
assign addr[38420]= -2040479063;
assign addr[38421]= -2015345591;
assign addr[38422]= -1987655498;
assign addr[38423]= -1957443913;
assign addr[38424]= -1924749160;
assign addr[38425]= -1889612716;
assign addr[38426]= -1852079154;
assign addr[38427]= -1812196087;
assign addr[38428]= -1770014111;
assign addr[38429]= -1725586737;
assign addr[38430]= -1678970324;
assign addr[38431]= -1630224009;
assign addr[38432]= -1579409630;
assign addr[38433]= -1526591649;
assign addr[38434]= -1471837070;
assign addr[38435]= -1415215352;
assign addr[38436]= -1356798326;
assign addr[38437]= -1296660098;
assign addr[38438]= -1234876957;
assign addr[38439]= -1171527280;
assign addr[38440]= -1106691431;
assign addr[38441]= -1040451659;
assign addr[38442]= -972891995;
assign addr[38443]= -904098143;
assign addr[38444]= -834157373;
assign addr[38445]= -763158411;
assign addr[38446]= -691191324;
assign addr[38447]= -618347408;
assign addr[38448]= -544719071;
assign addr[38449]= -470399716;
assign addr[38450]= -395483624;
assign addr[38451]= -320065829;
assign addr[38452]= -244242007;
assign addr[38453]= -168108346;
assign addr[38454]= -91761426;
assign addr[38455]= -15298099;
assign addr[38456]= 61184634;
assign addr[38457]= 137589750;
assign addr[38458]= 213820322;
assign addr[38459]= 289779648;
assign addr[38460]= 365371365;
assign addr[38461]= 440499581;
assign addr[38462]= 515068990;
assign addr[38463]= 588984994;
assign addr[38464]= 662153826;
assign addr[38465]= 734482665;
assign addr[38466]= 805879757;
assign addr[38467]= 876254528;
assign addr[38468]= 945517704;
assign addr[38469]= 1013581418;
assign addr[38470]= 1080359326;
assign addr[38471]= 1145766716;
assign addr[38472]= 1209720613;
assign addr[38473]= 1272139887;
assign addr[38474]= 1332945355;
assign addr[38475]= 1392059879;
assign addr[38476]= 1449408469;
assign addr[38477]= 1504918373;
assign addr[38478]= 1558519173;
assign addr[38479]= 1610142873;
assign addr[38480]= 1659723983;
assign addr[38481]= 1707199606;
assign addr[38482]= 1752509516;
assign addr[38483]= 1795596234;
assign addr[38484]= 1836405100;
assign addr[38485]= 1874884346;
assign addr[38486]= 1910985158;
assign addr[38487]= 1944661739;
assign addr[38488]= 1975871368;
assign addr[38489]= 2004574453;
assign addr[38490]= 2030734582;
assign addr[38491]= 2054318569;
assign addr[38492]= 2075296495;
assign addr[38493]= 2093641749;
assign addr[38494]= 2109331059;
assign addr[38495]= 2122344521;
assign addr[38496]= 2132665626;
assign addr[38497]= 2140281282;
assign addr[38498]= 2145181827;
assign addr[38499]= 2147361045;
assign addr[38500]= 2146816171;
assign addr[38501]= 2143547897;
assign addr[38502]= 2137560369;
assign addr[38503]= 2128861181;
assign addr[38504]= 2117461370;
assign addr[38505]= 2103375398;
assign addr[38506]= 2086621133;
assign addr[38507]= 2067219829;
assign addr[38508]= 2045196100;
assign addr[38509]= 2020577882;
assign addr[38510]= 1993396407;
assign addr[38511]= 1963686155;
assign addr[38512]= 1931484818;
assign addr[38513]= 1896833245;
assign addr[38514]= 1859775393;
assign addr[38515]= 1820358275;
assign addr[38516]= 1778631892;
assign addr[38517]= 1734649179;
assign addr[38518]= 1688465931;
assign addr[38519]= 1640140734;
assign addr[38520]= 1589734894;
assign addr[38521]= 1537312353;
assign addr[38522]= 1482939614;
assign addr[38523]= 1426685652;
assign addr[38524]= 1368621831;
assign addr[38525]= 1308821808;
assign addr[38526]= 1247361445;
assign addr[38527]= 1184318708;
assign addr[38528]= 1119773573;
assign addr[38529]= 1053807919;
assign addr[38530]= 986505429;
assign addr[38531]= 917951481;
assign addr[38532]= 848233042;
assign addr[38533]= 777438554;
assign addr[38534]= 705657826;
assign addr[38535]= 632981917;
assign addr[38536]= 559503022;
assign addr[38537]= 485314355;
assign addr[38538]= 410510029;
assign addr[38539]= 335184940;
assign addr[38540]= 259434643;
assign addr[38541]= 183355234;
assign addr[38542]= 107043224;
assign addr[38543]= 30595422;
assign addr[38544]= -45891193;
assign addr[38545]= -122319591;
assign addr[38546]= -198592817;
assign addr[38547]= -274614114;
assign addr[38548]= -350287041;
assign addr[38549]= -425515602;
assign addr[38550]= -500204365;
assign addr[38551]= -574258580;
assign addr[38552]= -647584304;
assign addr[38553]= -720088517;
assign addr[38554]= -791679244;
assign addr[38555]= -862265664;
assign addr[38556]= -931758235;
assign addr[38557]= -1000068799;
assign addr[38558]= -1067110699;
assign addr[38559]= -1132798888;
assign addr[38560]= -1197050035;
assign addr[38561]= -1259782632;
assign addr[38562]= -1320917099;
assign addr[38563]= -1380375881;
assign addr[38564]= -1438083551;
assign addr[38565]= -1493966902;
assign addr[38566]= -1547955041;
assign addr[38567]= -1599979481;
assign addr[38568]= -1649974225;
assign addr[38569]= -1697875851;
assign addr[38570]= -1743623590;
assign addr[38571]= -1787159411;
assign addr[38572]= -1828428082;
assign addr[38573]= -1867377253;
assign addr[38574]= -1903957513;
assign addr[38575]= -1938122457;
assign addr[38576]= -1969828744;
assign addr[38577]= -1999036154;
assign addr[38578]= -2025707632;
assign addr[38579]= -2049809346;
assign addr[38580]= -2071310720;
assign addr[38581]= -2090184478;
assign addr[38582]= -2106406677;
assign addr[38583]= -2119956737;
assign addr[38584]= -2130817471;
assign addr[38585]= -2138975100;
assign addr[38586]= -2144419275;
assign addr[38587]= -2147143090;
assign addr[38588]= -2147143090;
assign addr[38589]= -2144419275;
assign addr[38590]= -2138975100;
assign addr[38591]= -2130817471;
assign addr[38592]= -2119956737;
assign addr[38593]= -2106406677;
assign addr[38594]= -2090184478;
assign addr[38595]= -2071310720;
assign addr[38596]= -2049809346;
assign addr[38597]= -2025707632;
assign addr[38598]= -1999036154;
assign addr[38599]= -1969828744;
assign addr[38600]= -1938122457;
assign addr[38601]= -1903957513;
assign addr[38602]= -1867377253;
assign addr[38603]= -1828428082;
assign addr[38604]= -1787159411;
assign addr[38605]= -1743623590;
assign addr[38606]= -1697875851;
assign addr[38607]= -1649974225;
assign addr[38608]= -1599979481;
assign addr[38609]= -1547955041;
assign addr[38610]= -1493966902;
assign addr[38611]= -1438083551;
assign addr[38612]= -1380375881;
assign addr[38613]= -1320917099;
assign addr[38614]= -1259782632;
assign addr[38615]= -1197050035;
assign addr[38616]= -1132798888;
assign addr[38617]= -1067110699;
assign addr[38618]= -1000068799;
assign addr[38619]= -931758235;
assign addr[38620]= -862265664;
assign addr[38621]= -791679244;
assign addr[38622]= -720088517;
assign addr[38623]= -647584304;
assign addr[38624]= -574258580;
assign addr[38625]= -500204365;
assign addr[38626]= -425515602;
assign addr[38627]= -350287041;
assign addr[38628]= -274614114;
assign addr[38629]= -198592817;
assign addr[38630]= -122319591;
assign addr[38631]= -45891193;
assign addr[38632]= 30595422;
assign addr[38633]= 107043224;
assign addr[38634]= 183355234;
assign addr[38635]= 259434643;
assign addr[38636]= 335184940;
assign addr[38637]= 410510029;
assign addr[38638]= 485314355;
assign addr[38639]= 559503022;
assign addr[38640]= 632981917;
assign addr[38641]= 705657826;
assign addr[38642]= 777438554;
assign addr[38643]= 848233042;
assign addr[38644]= 917951481;
assign addr[38645]= 986505429;
assign addr[38646]= 1053807919;
assign addr[38647]= 1119773573;
assign addr[38648]= 1184318708;
assign addr[38649]= 1247361445;
assign addr[38650]= 1308821808;
assign addr[38651]= 1368621831;
assign addr[38652]= 1426685652;
assign addr[38653]= 1482939614;
assign addr[38654]= 1537312353;
assign addr[38655]= 1589734894;
assign addr[38656]= 1640140734;
assign addr[38657]= 1688465931;
assign addr[38658]= 1734649179;
assign addr[38659]= 1778631892;
assign addr[38660]= 1820358275;
assign addr[38661]= 1859775393;
assign addr[38662]= 1896833245;
assign addr[38663]= 1931484818;
assign addr[38664]= 1963686155;
assign addr[38665]= 1993396407;
assign addr[38666]= 2020577882;
assign addr[38667]= 2045196100;
assign addr[38668]= 2067219829;
assign addr[38669]= 2086621133;
assign addr[38670]= 2103375398;
assign addr[38671]= 2117461370;
assign addr[38672]= 2128861181;
assign addr[38673]= 2137560369;
assign addr[38674]= 2143547897;
assign addr[38675]= 2146816171;
assign addr[38676]= 2147361045;
assign addr[38677]= 2145181827;
assign addr[38678]= 2140281282;
assign addr[38679]= 2132665626;
assign addr[38680]= 2122344521;
assign addr[38681]= 2109331059;
assign addr[38682]= 2093641749;
assign addr[38683]= 2075296495;
assign addr[38684]= 2054318569;
assign addr[38685]= 2030734582;
assign addr[38686]= 2004574453;
assign addr[38687]= 1975871368;
assign addr[38688]= 1944661739;
assign addr[38689]= 1910985158;
assign addr[38690]= 1874884346;
assign addr[38691]= 1836405100;
assign addr[38692]= 1795596234;
assign addr[38693]= 1752509516;
assign addr[38694]= 1707199606;
assign addr[38695]= 1659723983;
assign addr[38696]= 1610142873;
assign addr[38697]= 1558519173;
assign addr[38698]= 1504918373;
assign addr[38699]= 1449408469;
assign addr[38700]= 1392059879;
assign addr[38701]= 1332945355;
assign addr[38702]= 1272139887;
assign addr[38703]= 1209720613;
assign addr[38704]= 1145766716;
assign addr[38705]= 1080359326;
assign addr[38706]= 1013581418;
assign addr[38707]= 945517704;
assign addr[38708]= 876254528;
assign addr[38709]= 805879757;
assign addr[38710]= 734482665;
assign addr[38711]= 662153826;
assign addr[38712]= 588984994;
assign addr[38713]= 515068990;
assign addr[38714]= 440499581;
assign addr[38715]= 365371365;
assign addr[38716]= 289779648;
assign addr[38717]= 213820322;
assign addr[38718]= 137589750;
assign addr[38719]= 61184634;
assign addr[38720]= -15298099;
assign addr[38721]= -91761426;
assign addr[38722]= -168108346;
assign addr[38723]= -244242007;
assign addr[38724]= -320065829;
assign addr[38725]= -395483624;
assign addr[38726]= -470399716;
assign addr[38727]= -544719071;
assign addr[38728]= -618347408;
assign addr[38729]= -691191324;
assign addr[38730]= -763158411;
assign addr[38731]= -834157373;
assign addr[38732]= -904098143;
assign addr[38733]= -972891995;
assign addr[38734]= -1040451659;
assign addr[38735]= -1106691431;
assign addr[38736]= -1171527280;
assign addr[38737]= -1234876957;
assign addr[38738]= -1296660098;
assign addr[38739]= -1356798326;
assign addr[38740]= -1415215352;
assign addr[38741]= -1471837070;
assign addr[38742]= -1526591649;
assign addr[38743]= -1579409630;
assign addr[38744]= -1630224009;
assign addr[38745]= -1678970324;
assign addr[38746]= -1725586737;
assign addr[38747]= -1770014111;
assign addr[38748]= -1812196087;
assign addr[38749]= -1852079154;
assign addr[38750]= -1889612716;
assign addr[38751]= -1924749160;
assign addr[38752]= -1957443913;
assign addr[38753]= -1987655498;
assign addr[38754]= -2015345591;
assign addr[38755]= -2040479063;
assign addr[38756]= -2063024031;
assign addr[38757]= -2082951896;
assign addr[38758]= -2100237377;
assign addr[38759]= -2114858546;
assign addr[38760]= -2126796855;
assign addr[38761]= -2136037160;
assign addr[38762]= -2142567738;
assign addr[38763]= -2146380306;
assign addr[38764]= -2147470025;
assign addr[38765]= -2145835515;
assign addr[38766]= -2141478848;
assign addr[38767]= -2134405552;
assign addr[38768]= -2124624598;
assign addr[38769]= -2112148396;
assign addr[38770]= -2096992772;
assign addr[38771]= -2079176953;
assign addr[38772]= -2058723538;
assign addr[38773]= -2035658475;
assign addr[38774]= -2010011024;
assign addr[38775]= -1981813720;
assign addr[38776]= -1951102334;
assign addr[38777]= -1917915825;
assign addr[38778]= -1882296293;
assign addr[38779]= -1844288924;
assign addr[38780]= -1803941934;
assign addr[38781]= -1761306505;
assign addr[38782]= -1716436725;
assign addr[38783]= -1669389513;
assign addr[38784]= -1620224553;
assign addr[38785]= -1569004214;
assign addr[38786]= -1515793473;
assign addr[38787]= -1460659832;
assign addr[38788]= -1403673233;
assign addr[38789]= -1344905966;
assign addr[38790]= -1284432584;
assign addr[38791]= -1222329801;
assign addr[38792]= -1158676398;
assign addr[38793]= -1093553126;
assign addr[38794]= -1027042599;
assign addr[38795]= -959229189;
assign addr[38796]= -890198924;
assign addr[38797]= -820039373;
assign addr[38798]= -748839539;
assign addr[38799]= -676689746;
assign addr[38800]= -603681519;
assign addr[38801]= -529907477;
assign addr[38802]= -455461206;
assign addr[38803]= -380437148;
assign addr[38804]= -304930476;
assign addr[38805]= -229036977;
assign addr[38806]= -152852926;
assign addr[38807]= -76474970;
assign addr[38808]= 0;
assign addr[38809]= 76474970;
assign addr[38810]= 152852926;
assign addr[38811]= 229036977;
assign addr[38812]= 304930476;
assign addr[38813]= 380437148;
assign addr[38814]= 455461206;
assign addr[38815]= 529907477;
assign addr[38816]= 603681519;
assign addr[38817]= 676689746;
assign addr[38818]= 748839539;
assign addr[38819]= 820039373;
assign addr[38820]= 890198924;
assign addr[38821]= 959229189;
assign addr[38822]= 1027042599;
assign addr[38823]= 1093553126;
assign addr[38824]= 1158676398;
assign addr[38825]= 1222329801;
assign addr[38826]= 1284432584;
assign addr[38827]= 1344905966;
assign addr[38828]= 1403673233;
assign addr[38829]= 1460659832;
assign addr[38830]= 1515793473;
assign addr[38831]= 1569004214;
assign addr[38832]= 1620224553;
assign addr[38833]= 1669389513;
assign addr[38834]= 1716436725;
assign addr[38835]= 1761306505;
assign addr[38836]= 1803941934;
assign addr[38837]= 1844288924;
assign addr[38838]= 1882296293;
assign addr[38839]= 1917915825;
assign addr[38840]= 1951102334;
assign addr[38841]= 1981813720;
assign addr[38842]= 2010011024;
assign addr[38843]= 2035658475;
assign addr[38844]= 2058723538;
assign addr[38845]= 2079176953;
assign addr[38846]= 2096992772;
assign addr[38847]= 2112148396;
assign addr[38848]= 2124624598;
assign addr[38849]= 2134405552;
assign addr[38850]= 2141478848;
assign addr[38851]= 2145835515;
assign addr[38852]= 2147470025;
assign addr[38853]= 2146380306;
assign addr[38854]= 2142567738;
assign addr[38855]= 2136037160;
assign addr[38856]= 2126796855;
assign addr[38857]= 2114858546;
assign addr[38858]= 2100237377;
assign addr[38859]= 2082951896;
assign addr[38860]= 2063024031;
assign addr[38861]= 2040479063;
assign addr[38862]= 2015345591;
assign addr[38863]= 1987655498;
assign addr[38864]= 1957443913;
assign addr[38865]= 1924749160;
assign addr[38866]= 1889612716;
assign addr[38867]= 1852079154;
assign addr[38868]= 1812196087;
assign addr[38869]= 1770014111;
assign addr[38870]= 1725586737;
assign addr[38871]= 1678970324;
assign addr[38872]= 1630224009;
assign addr[38873]= 1579409630;
assign addr[38874]= 1526591649;
assign addr[38875]= 1471837070;
assign addr[38876]= 1415215352;
assign addr[38877]= 1356798326;
assign addr[38878]= 1296660098;
assign addr[38879]= 1234876957;
assign addr[38880]= 1171527280;
assign addr[38881]= 1106691431;
assign addr[38882]= 1040451659;
assign addr[38883]= 972891995;
assign addr[38884]= 904098143;
assign addr[38885]= 834157373;
assign addr[38886]= 763158411;
assign addr[38887]= 691191324;
assign addr[38888]= 618347408;
assign addr[38889]= 544719071;
assign addr[38890]= 470399716;
assign addr[38891]= 395483624;
assign addr[38892]= 320065829;
assign addr[38893]= 244242007;
assign addr[38894]= 168108346;
assign addr[38895]= 91761426;
assign addr[38896]= 15298099;
assign addr[38897]= -61184634;
assign addr[38898]= -137589750;
assign addr[38899]= -213820322;
assign addr[38900]= -289779648;
assign addr[38901]= -365371365;
assign addr[38902]= -440499581;
assign addr[38903]= -515068990;
assign addr[38904]= -588984994;
assign addr[38905]= -662153826;
assign addr[38906]= -734482665;
assign addr[38907]= -805879757;
assign addr[38908]= -876254528;
assign addr[38909]= -945517704;
assign addr[38910]= -1013581418;
assign addr[38911]= -1080359326;
assign addr[38912]= -1145766716;
assign addr[38913]= -1209720613;
assign addr[38914]= -1272139887;
assign addr[38915]= -1332945355;
assign addr[38916]= -1392059879;
assign addr[38917]= -1449408469;
assign addr[38918]= -1504918373;
assign addr[38919]= -1558519173;
assign addr[38920]= -1610142873;
assign addr[38921]= -1659723983;
assign addr[38922]= -1707199606;
assign addr[38923]= -1752509516;
assign addr[38924]= -1795596234;
assign addr[38925]= -1836405100;
assign addr[38926]= -1874884346;
assign addr[38927]= -1910985158;
assign addr[38928]= -1944661739;
assign addr[38929]= -1975871368;
assign addr[38930]= -2004574453;
assign addr[38931]= -2030734582;
assign addr[38932]= -2054318569;
assign addr[38933]= -2075296495;
assign addr[38934]= -2093641749;
assign addr[38935]= -2109331059;
assign addr[38936]= -2122344521;
assign addr[38937]= -2132665626;
assign addr[38938]= -2140281282;
assign addr[38939]= -2145181827;
assign addr[38940]= -2147361045;
assign addr[38941]= -2146816171;
assign addr[38942]= -2143547897;
assign addr[38943]= -2137560369;
assign addr[38944]= -2128861181;
assign addr[38945]= -2117461370;
assign addr[38946]= -2103375398;
assign addr[38947]= -2086621133;
assign addr[38948]= -2067219829;
assign addr[38949]= -2045196100;
assign addr[38950]= -2020577882;
assign addr[38951]= -1993396407;
assign addr[38952]= -1963686155;
assign addr[38953]= -1931484818;
assign addr[38954]= -1896833245;
assign addr[38955]= -1859775393;
assign addr[38956]= -1820358275;
assign addr[38957]= -1778631892;
assign addr[38958]= -1734649179;
assign addr[38959]= -1688465931;
assign addr[38960]= -1640140734;
assign addr[38961]= -1589734894;
assign addr[38962]= -1537312353;
assign addr[38963]= -1482939614;
assign addr[38964]= -1426685652;
assign addr[38965]= -1368621831;
assign addr[38966]= -1308821808;
assign addr[38967]= -1247361445;
assign addr[38968]= -1184318708;
assign addr[38969]= -1119773573;
assign addr[38970]= -1053807919;
assign addr[38971]= -986505429;
assign addr[38972]= -917951481;
assign addr[38973]= -848233042;
assign addr[38974]= -777438554;
assign addr[38975]= -705657826;
assign addr[38976]= -632981917;
assign addr[38977]= -559503022;
assign addr[38978]= -485314355;
assign addr[38979]= -410510029;
assign addr[38980]= -335184940;
assign addr[38981]= -259434643;
assign addr[38982]= -183355234;
assign addr[38983]= -107043224;
assign addr[38984]= -30595422;
assign addr[38985]= 45891193;
assign addr[38986]= 122319591;
assign addr[38987]= 198592817;
assign addr[38988]= 274614114;
assign addr[38989]= 350287041;
assign addr[38990]= 425515602;
assign addr[38991]= 500204365;
assign addr[38992]= 574258580;
assign addr[38993]= 647584304;
assign addr[38994]= 720088517;
assign addr[38995]= 791679244;
assign addr[38996]= 862265664;
assign addr[38997]= 931758235;
assign addr[38998]= 1000068799;
assign addr[38999]= 1067110699;
assign addr[39000]= 1132798888;
assign addr[39001]= 1197050035;
assign addr[39002]= 1259782632;
assign addr[39003]= 1320917099;
assign addr[39004]= 1380375881;
assign addr[39005]= 1438083551;
assign addr[39006]= 1493966902;
assign addr[39007]= 1547955041;
assign addr[39008]= 1599979481;
assign addr[39009]= 1649974225;
assign addr[39010]= 1697875851;
assign addr[39011]= 1743623590;
assign addr[39012]= 1787159411;
assign addr[39013]= 1828428082;
assign addr[39014]= 1867377253;
assign addr[39015]= 1903957513;
assign addr[39016]= 1938122457;
assign addr[39017]= 1969828744;
assign addr[39018]= 1999036154;
assign addr[39019]= 2025707632;
assign addr[39020]= 2049809346;
assign addr[39021]= 2071310720;
assign addr[39022]= 2090184478;
assign addr[39023]= 2106406677;
assign addr[39024]= 2119956737;
assign addr[39025]= 2130817471;
assign addr[39026]= 2138975100;
assign addr[39027]= 2144419275;
assign addr[39028]= 2147143090;
assign addr[39029]= 2147143090;
assign addr[39030]= 2144419275;
assign addr[39031]= 2138975100;
assign addr[39032]= 2130817471;
assign addr[39033]= 2119956737;
assign addr[39034]= 2106406677;
assign addr[39035]= 2090184478;
assign addr[39036]= 2071310720;
assign addr[39037]= 2049809346;
assign addr[39038]= 2025707632;
assign addr[39039]= 1999036154;
assign addr[39040]= 1969828744;
assign addr[39041]= 1938122457;
assign addr[39042]= 1903957513;
assign addr[39043]= 1867377253;
assign addr[39044]= 1828428082;
assign addr[39045]= 1787159411;
assign addr[39046]= 1743623590;
assign addr[39047]= 1697875851;
assign addr[39048]= 1649974225;
assign addr[39049]= 1599979481;
assign addr[39050]= 1547955041;
assign addr[39051]= 1493966902;
assign addr[39052]= 1438083551;
assign addr[39053]= 1380375881;
assign addr[39054]= 1320917099;
assign addr[39055]= 1259782632;
assign addr[39056]= 1197050035;
assign addr[39057]= 1132798888;
assign addr[39058]= 1067110699;
assign addr[39059]= 1000068799;
assign addr[39060]= 931758235;
assign addr[39061]= 862265664;
assign addr[39062]= 791679244;
assign addr[39063]= 720088517;
assign addr[39064]= 647584304;
assign addr[39065]= 574258580;
assign addr[39066]= 500204365;
assign addr[39067]= 425515602;
assign addr[39068]= 350287041;
assign addr[39069]= 274614114;
assign addr[39070]= 198592817;
assign addr[39071]= 122319591;
assign addr[39072]= 45891193;
assign addr[39073]= -30595422;
assign addr[39074]= -107043224;
assign addr[39075]= -183355234;
assign addr[39076]= -259434643;
assign addr[39077]= -335184940;
assign addr[39078]= -410510029;
assign addr[39079]= -485314355;
assign addr[39080]= -559503022;
assign addr[39081]= -632981917;
assign addr[39082]= -705657826;
assign addr[39083]= -777438554;
assign addr[39084]= -848233042;
assign addr[39085]= -917951481;
assign addr[39086]= -986505429;
assign addr[39087]= -1053807919;
assign addr[39088]= -1119773573;
assign addr[39089]= -1184318708;
assign addr[39090]= -1247361445;
assign addr[39091]= -1308821808;
assign addr[39092]= -1368621831;
assign addr[39093]= -1426685652;
assign addr[39094]= -1482939614;
assign addr[39095]= -1537312353;
assign addr[39096]= -1589734894;
assign addr[39097]= -1640140734;
assign addr[39098]= -1688465931;
assign addr[39099]= -1734649179;
assign addr[39100]= -1778631892;
assign addr[39101]= -1820358275;
assign addr[39102]= -1859775393;
assign addr[39103]= -1896833245;
assign addr[39104]= -1931484818;
assign addr[39105]= -1963686155;
assign addr[39106]= -1993396407;
assign addr[39107]= -2020577882;
assign addr[39108]= -2045196100;
assign addr[39109]= -2067219829;
assign addr[39110]= -2086621133;
assign addr[39111]= -2103375398;
assign addr[39112]= -2117461370;
assign addr[39113]= -2128861181;
assign addr[39114]= -2137560369;
assign addr[39115]= -2143547897;
assign addr[39116]= -2146816171;
assign addr[39117]= -2147361045;
assign addr[39118]= -2145181827;
assign addr[39119]= -2140281282;
assign addr[39120]= -2132665626;
assign addr[39121]= -2122344521;
assign addr[39122]= -2109331059;
assign addr[39123]= -2093641749;
assign addr[39124]= -2075296495;
assign addr[39125]= -2054318569;
assign addr[39126]= -2030734582;
assign addr[39127]= -2004574453;
assign addr[39128]= -1975871368;
assign addr[39129]= -1944661739;
assign addr[39130]= -1910985158;
assign addr[39131]= -1874884346;
assign addr[39132]= -1836405100;
assign addr[39133]= -1795596234;
assign addr[39134]= -1752509516;
assign addr[39135]= -1707199606;
assign addr[39136]= -1659723983;
assign addr[39137]= -1610142873;
assign addr[39138]= -1558519173;
assign addr[39139]= -1504918373;
assign addr[39140]= -1449408469;
assign addr[39141]= -1392059879;
assign addr[39142]= -1332945355;
assign addr[39143]= -1272139887;
assign addr[39144]= -1209720613;
assign addr[39145]= -1145766716;
assign addr[39146]= -1080359326;
assign addr[39147]= -1013581418;
assign addr[39148]= -945517704;
assign addr[39149]= -876254528;
assign addr[39150]= -805879757;
assign addr[39151]= -734482665;
assign addr[39152]= -662153826;
assign addr[39153]= -588984994;
assign addr[39154]= -515068990;
assign addr[39155]= -440499581;
assign addr[39156]= -365371365;
assign addr[39157]= -289779648;
assign addr[39158]= -213820322;
assign addr[39159]= -137589750;
assign addr[39160]= -61184634;
assign addr[39161]= 15298099;
assign addr[39162]= 91761426;
assign addr[39163]= 168108346;
assign addr[39164]= 244242007;
assign addr[39165]= 320065829;
assign addr[39166]= 395483624;
assign addr[39167]= 470399716;
assign addr[39168]= 544719071;
assign addr[39169]= 618347408;
assign addr[39170]= 691191324;
assign addr[39171]= 763158411;
assign addr[39172]= 834157373;
assign addr[39173]= 904098143;
assign addr[39174]= 972891995;
assign addr[39175]= 1040451659;
assign addr[39176]= 1106691431;
assign addr[39177]= 1171527280;
assign addr[39178]= 1234876957;
assign addr[39179]= 1296660098;
assign addr[39180]= 1356798326;
assign addr[39181]= 1415215352;
assign addr[39182]= 1471837070;
assign addr[39183]= 1526591649;
assign addr[39184]= 1579409630;
assign addr[39185]= 1630224009;
assign addr[39186]= 1678970324;
assign addr[39187]= 1725586737;
assign addr[39188]= 1770014111;
assign addr[39189]= 1812196087;
assign addr[39190]= 1852079154;
assign addr[39191]= 1889612716;
assign addr[39192]= 1924749160;
assign addr[39193]= 1957443913;
assign addr[39194]= 1987655498;
assign addr[39195]= 2015345591;
assign addr[39196]= 2040479063;
assign addr[39197]= 2063024031;
assign addr[39198]= 2082951896;
assign addr[39199]= 2100237377;
assign addr[39200]= 2114858546;
assign addr[39201]= 2126796855;
assign addr[39202]= 2136037160;
assign addr[39203]= 2142567738;
assign addr[39204]= 2146380306;
assign addr[39205]= 2147470025;
assign addr[39206]= 2145835515;
assign addr[39207]= 2141478848;
assign addr[39208]= 2134405552;
assign addr[39209]= 2124624598;
assign addr[39210]= 2112148396;
assign addr[39211]= 2096992772;
assign addr[39212]= 2079176953;
assign addr[39213]= 2058723538;
assign addr[39214]= 2035658475;
assign addr[39215]= 2010011024;
assign addr[39216]= 1981813720;
assign addr[39217]= 1951102334;
assign addr[39218]= 1917915825;
assign addr[39219]= 1882296293;
assign addr[39220]= 1844288924;
assign addr[39221]= 1803941934;
assign addr[39222]= 1761306505;
assign addr[39223]= 1716436725;
assign addr[39224]= 1669389513;
assign addr[39225]= 1620224553;
assign addr[39226]= 1569004214;
assign addr[39227]= 1515793473;
assign addr[39228]= 1460659832;
assign addr[39229]= 1403673233;
assign addr[39230]= 1344905966;
assign addr[39231]= 1284432584;
assign addr[39232]= 1222329801;
assign addr[39233]= 1158676398;
assign addr[39234]= 1093553126;
assign addr[39235]= 1027042599;
assign addr[39236]= 959229189;
assign addr[39237]= 890198924;
assign addr[39238]= 820039373;
assign addr[39239]= 748839539;
assign addr[39240]= 676689746;
assign addr[39241]= 603681519;
assign addr[39242]= 529907477;
assign addr[39243]= 455461206;
assign addr[39244]= 380437148;
assign addr[39245]= 304930476;
assign addr[39246]= 229036977;
assign addr[39247]= 152852926;
assign addr[39248]= 76474970;
assign addr[39249]= 0;
assign addr[39250]= -76474970;
assign addr[39251]= -152852926;
assign addr[39252]= -229036977;
assign addr[39253]= -304930476;
assign addr[39254]= -380437148;
assign addr[39255]= -455461206;
assign addr[39256]= -529907477;
assign addr[39257]= -603681519;
assign addr[39258]= -676689746;
assign addr[39259]= -748839539;
assign addr[39260]= -820039373;
assign addr[39261]= -890198924;
assign addr[39262]= -959229189;
assign addr[39263]= -1027042599;
assign addr[39264]= -1093553126;
assign addr[39265]= -1158676398;
assign addr[39266]= -1222329801;
assign addr[39267]= -1284432584;
assign addr[39268]= -1344905966;
assign addr[39269]= -1403673233;
assign addr[39270]= -1460659832;
assign addr[39271]= -1515793473;
assign addr[39272]= -1569004214;
assign addr[39273]= -1620224553;
assign addr[39274]= -1669389513;
assign addr[39275]= -1716436725;
assign addr[39276]= -1761306505;
assign addr[39277]= -1803941934;
assign addr[39278]= -1844288924;
assign addr[39279]= -1882296293;
assign addr[39280]= -1917915825;
assign addr[39281]= -1951102334;
assign addr[39282]= -1981813720;
assign addr[39283]= -2010011024;
assign addr[39284]= -2035658475;
assign addr[39285]= -2058723538;
assign addr[39286]= -2079176953;
assign addr[39287]= -2096992772;
assign addr[39288]= -2112148396;
assign addr[39289]= -2124624598;
assign addr[39290]= -2134405552;
assign addr[39291]= -2141478848;
assign addr[39292]= -2145835515;
assign addr[39293]= -2147470025;
assign addr[39294]= -2146380306;
assign addr[39295]= -2142567738;
assign addr[39296]= -2136037160;
assign addr[39297]= -2126796855;
assign addr[39298]= -2114858546;
assign addr[39299]= -2100237377;
assign addr[39300]= -2082951896;
assign addr[39301]= -2063024031;
assign addr[39302]= -2040479063;
assign addr[39303]= -2015345591;
assign addr[39304]= -1987655498;
assign addr[39305]= -1957443913;
assign addr[39306]= -1924749160;
assign addr[39307]= -1889612716;
assign addr[39308]= -1852079154;
assign addr[39309]= -1812196087;
assign addr[39310]= -1770014111;
assign addr[39311]= -1725586737;
assign addr[39312]= -1678970324;
assign addr[39313]= -1630224009;
assign addr[39314]= -1579409630;
assign addr[39315]= -1526591649;
assign addr[39316]= -1471837070;
assign addr[39317]= -1415215352;
assign addr[39318]= -1356798326;
assign addr[39319]= -1296660098;
assign addr[39320]= -1234876957;
assign addr[39321]= -1171527280;
assign addr[39322]= -1106691431;
assign addr[39323]= -1040451659;
assign addr[39324]= -972891995;
assign addr[39325]= -904098143;
assign addr[39326]= -834157373;
assign addr[39327]= -763158411;
assign addr[39328]= -691191324;
assign addr[39329]= -618347408;
assign addr[39330]= -544719071;
assign addr[39331]= -470399716;
assign addr[39332]= -395483624;
assign addr[39333]= -320065829;
assign addr[39334]= -244242007;
assign addr[39335]= -168108346;
assign addr[39336]= -91761426;
assign addr[39337]= -15298099;
assign addr[39338]= 61184634;
assign addr[39339]= 137589750;
assign addr[39340]= 213820322;
assign addr[39341]= 289779648;
assign addr[39342]= 365371365;
assign addr[39343]= 440499581;
assign addr[39344]= 515068990;
assign addr[39345]= 588984994;
assign addr[39346]= 662153826;
assign addr[39347]= 734482665;
assign addr[39348]= 805879757;
assign addr[39349]= 876254528;
assign addr[39350]= 945517704;
assign addr[39351]= 1013581418;
assign addr[39352]= 1080359326;
assign addr[39353]= 1145766716;
assign addr[39354]= 1209720613;
assign addr[39355]= 1272139887;
assign addr[39356]= 1332945355;
assign addr[39357]= 1392059879;
assign addr[39358]= 1449408469;
assign addr[39359]= 1504918373;
assign addr[39360]= 1558519173;
assign addr[39361]= 1610142873;
assign addr[39362]= 1659723983;
assign addr[39363]= 1707199606;
assign addr[39364]= 1752509516;
assign addr[39365]= 1795596234;
assign addr[39366]= 1836405100;
assign addr[39367]= 1874884346;
assign addr[39368]= 1910985158;
assign addr[39369]= 1944661739;
assign addr[39370]= 1975871368;
assign addr[39371]= 2004574453;
assign addr[39372]= 2030734582;
assign addr[39373]= 2054318569;
assign addr[39374]= 2075296495;
assign addr[39375]= 2093641749;
assign addr[39376]= 2109331059;
assign addr[39377]= 2122344521;
assign addr[39378]= 2132665626;
assign addr[39379]= 2140281282;
assign addr[39380]= 2145181827;
assign addr[39381]= 2147361045;
assign addr[39382]= 2146816171;
assign addr[39383]= 2143547897;
assign addr[39384]= 2137560369;
assign addr[39385]= 2128861181;
assign addr[39386]= 2117461370;
assign addr[39387]= 2103375398;
assign addr[39388]= 2086621133;
assign addr[39389]= 2067219829;
assign addr[39390]= 2045196100;
assign addr[39391]= 2020577882;
assign addr[39392]= 1993396407;
assign addr[39393]= 1963686155;
assign addr[39394]= 1931484818;
assign addr[39395]= 1896833245;
assign addr[39396]= 1859775393;
assign addr[39397]= 1820358275;
assign addr[39398]= 1778631892;
assign addr[39399]= 1734649179;
assign addr[39400]= 1688465931;
assign addr[39401]= 1640140734;
assign addr[39402]= 1589734894;
assign addr[39403]= 1537312353;
assign addr[39404]= 1482939614;
assign addr[39405]= 1426685652;
assign addr[39406]= 1368621831;
assign addr[39407]= 1308821808;
assign addr[39408]= 1247361445;
assign addr[39409]= 1184318708;
assign addr[39410]= 1119773573;
assign addr[39411]= 1053807919;
assign addr[39412]= 986505429;
assign addr[39413]= 917951481;
assign addr[39414]= 848233042;
assign addr[39415]= 777438554;
assign addr[39416]= 705657826;
assign addr[39417]= 632981917;
assign addr[39418]= 559503022;
assign addr[39419]= 485314355;
assign addr[39420]= 410510029;
assign addr[39421]= 335184940;
assign addr[39422]= 259434643;
assign addr[39423]= 183355234;
assign addr[39424]= 107043224;
assign addr[39425]= 30595422;
assign addr[39426]= -45891193;
assign addr[39427]= -122319591;
assign addr[39428]= -198592817;
assign addr[39429]= -274614114;
assign addr[39430]= -350287041;
assign addr[39431]= -425515602;
assign addr[39432]= -500204365;
assign addr[39433]= -574258580;
assign addr[39434]= -647584304;
assign addr[39435]= -720088517;
assign addr[39436]= -791679244;
assign addr[39437]= -862265664;
assign addr[39438]= -931758235;
assign addr[39439]= -1000068799;
assign addr[39440]= -1067110699;
assign addr[39441]= -1132798888;
assign addr[39442]= -1197050035;
assign addr[39443]= -1259782632;
assign addr[39444]= -1320917099;
assign addr[39445]= -1380375881;
assign addr[39446]= -1438083551;
assign addr[39447]= -1493966902;
assign addr[39448]= -1547955041;
assign addr[39449]= -1599979481;
assign addr[39450]= -1649974225;
assign addr[39451]= -1697875851;
assign addr[39452]= -1743623590;
assign addr[39453]= -1787159411;
assign addr[39454]= -1828428082;
assign addr[39455]= -1867377253;
assign addr[39456]= -1903957513;
assign addr[39457]= -1938122457;
assign addr[39458]= -1969828744;
assign addr[39459]= -1999036154;
assign addr[39460]= -2025707632;
assign addr[39461]= -2049809346;
assign addr[39462]= -2071310720;
assign addr[39463]= -2090184478;
assign addr[39464]= -2106406677;
assign addr[39465]= -2119956737;
assign addr[39466]= -2130817471;
assign addr[39467]= -2138975100;
assign addr[39468]= -2144419275;
assign addr[39469]= -2147143090;
assign addr[39470]= -2147143090;
assign addr[39471]= -2144419275;
assign addr[39472]= -2138975100;
assign addr[39473]= -2130817471;
assign addr[39474]= -2119956737;
assign addr[39475]= -2106406677;
assign addr[39476]= -2090184478;
assign addr[39477]= -2071310720;
assign addr[39478]= -2049809346;
assign addr[39479]= -2025707632;
assign addr[39480]= -1999036154;
assign addr[39481]= -1969828744;
assign addr[39482]= -1938122457;
assign addr[39483]= -1903957513;
assign addr[39484]= -1867377253;
assign addr[39485]= -1828428082;
assign addr[39486]= -1787159411;
assign addr[39487]= -1743623590;
assign addr[39488]= -1697875851;
assign addr[39489]= -1649974225;
assign addr[39490]= -1599979481;
assign addr[39491]= -1547955041;
assign addr[39492]= -1493966902;
assign addr[39493]= -1438083551;
assign addr[39494]= -1380375881;
assign addr[39495]= -1320917099;
assign addr[39496]= -1259782632;
assign addr[39497]= -1197050035;
assign addr[39498]= -1132798888;
assign addr[39499]= -1067110699;
assign addr[39500]= -1000068799;
assign addr[39501]= -931758235;
assign addr[39502]= -862265664;
assign addr[39503]= -791679244;
assign addr[39504]= -720088517;
assign addr[39505]= -647584304;
assign addr[39506]= -574258580;
assign addr[39507]= -500204365;
assign addr[39508]= -425515602;
assign addr[39509]= -350287041;
assign addr[39510]= -274614114;
assign addr[39511]= -198592817;
assign addr[39512]= -122319591;
assign addr[39513]= -45891193;
assign addr[39514]= 30595422;
assign addr[39515]= 107043224;
assign addr[39516]= 183355234;
assign addr[39517]= 259434643;
assign addr[39518]= 335184940;
assign addr[39519]= 410510029;
assign addr[39520]= 485314355;
assign addr[39521]= 559503022;
assign addr[39522]= 632981917;
assign addr[39523]= 705657826;
assign addr[39524]= 777438554;
assign addr[39525]= 848233042;
assign addr[39526]= 917951481;
assign addr[39527]= 986505429;
assign addr[39528]= 1053807919;
assign addr[39529]= 1119773573;
assign addr[39530]= 1184318708;
assign addr[39531]= 1247361445;
assign addr[39532]= 1308821808;
assign addr[39533]= 1368621831;
assign addr[39534]= 1426685652;
assign addr[39535]= 1482939614;
assign addr[39536]= 1537312353;
assign addr[39537]= 1589734894;
assign addr[39538]= 1640140734;
assign addr[39539]= 1688465931;
assign addr[39540]= 1734649179;
assign addr[39541]= 1778631892;
assign addr[39542]= 1820358275;
assign addr[39543]= 1859775393;
assign addr[39544]= 1896833245;
assign addr[39545]= 1931484818;
assign addr[39546]= 1963686155;
assign addr[39547]= 1993396407;
assign addr[39548]= 2020577882;
assign addr[39549]= 2045196100;
assign addr[39550]= 2067219829;
assign addr[39551]= 2086621133;
assign addr[39552]= 2103375398;
assign addr[39553]= 2117461370;
assign addr[39554]= 2128861181;
assign addr[39555]= 2137560369;
assign addr[39556]= 2143547897;
assign addr[39557]= 2146816171;
assign addr[39558]= 2147361045;
assign addr[39559]= 2145181827;
assign addr[39560]= 2140281282;
assign addr[39561]= 2132665626;
assign addr[39562]= 2122344521;
assign addr[39563]= 2109331059;
assign addr[39564]= 2093641749;
assign addr[39565]= 2075296495;
assign addr[39566]= 2054318569;
assign addr[39567]= 2030734582;
assign addr[39568]= 2004574453;
assign addr[39569]= 1975871368;
assign addr[39570]= 1944661739;
assign addr[39571]= 1910985158;
assign addr[39572]= 1874884346;
assign addr[39573]= 1836405100;
assign addr[39574]= 1795596234;
assign addr[39575]= 1752509516;
assign addr[39576]= 1707199606;
assign addr[39577]= 1659723983;
assign addr[39578]= 1610142873;
assign addr[39579]= 1558519173;
assign addr[39580]= 1504918373;
assign addr[39581]= 1449408469;
assign addr[39582]= 1392059879;
assign addr[39583]= 1332945355;
assign addr[39584]= 1272139887;
assign addr[39585]= 1209720613;
assign addr[39586]= 1145766716;
assign addr[39587]= 1080359326;
assign addr[39588]= 1013581418;
assign addr[39589]= 945517704;
assign addr[39590]= 876254528;
assign addr[39591]= 805879757;
assign addr[39592]= 734482665;
assign addr[39593]= 662153826;
assign addr[39594]= 588984994;
assign addr[39595]= 515068990;
assign addr[39596]= 440499581;
assign addr[39597]= 365371365;
assign addr[39598]= 289779648;
assign addr[39599]= 213820322;
assign addr[39600]= 137589750;
assign addr[39601]= 61184634;
assign addr[39602]= -15298099;
assign addr[39603]= -91761426;
assign addr[39604]= -168108346;
assign addr[39605]= -244242007;
assign addr[39606]= -320065829;
assign addr[39607]= -395483624;
assign addr[39608]= -470399716;
assign addr[39609]= -544719071;
assign addr[39610]= -618347408;
assign addr[39611]= -691191324;
assign addr[39612]= -763158411;
assign addr[39613]= -834157373;
assign addr[39614]= -904098143;
assign addr[39615]= -972891995;
assign addr[39616]= -1040451659;
assign addr[39617]= -1106691431;
assign addr[39618]= -1171527280;
assign addr[39619]= -1234876957;
assign addr[39620]= -1296660098;
assign addr[39621]= -1356798326;
assign addr[39622]= -1415215352;
assign addr[39623]= -1471837070;
assign addr[39624]= -1526591649;
assign addr[39625]= -1579409630;
assign addr[39626]= -1630224009;
assign addr[39627]= -1678970324;
assign addr[39628]= -1725586737;
assign addr[39629]= -1770014111;
assign addr[39630]= -1812196087;
assign addr[39631]= -1852079154;
assign addr[39632]= -1889612716;
assign addr[39633]= -1924749160;
assign addr[39634]= -1957443913;
assign addr[39635]= -1987655498;
assign addr[39636]= -2015345591;
assign addr[39637]= -2040479063;
assign addr[39638]= -2063024031;
assign addr[39639]= -2082951896;
assign addr[39640]= -2100237377;
assign addr[39641]= -2114858546;
assign addr[39642]= -2126796855;
assign addr[39643]= -2136037160;
assign addr[39644]= -2142567738;
assign addr[39645]= -2146380306;
assign addr[39646]= -2147470025;
assign addr[39647]= -2145835515;
assign addr[39648]= -2141478848;
assign addr[39649]= -2134405552;
assign addr[39650]= -2124624598;
assign addr[39651]= -2112148396;
assign addr[39652]= -2096992772;
assign addr[39653]= -2079176953;
assign addr[39654]= -2058723538;
assign addr[39655]= -2035658475;
assign addr[39656]= -2010011024;
assign addr[39657]= -1981813720;
assign addr[39658]= -1951102334;
assign addr[39659]= -1917915825;
assign addr[39660]= -1882296293;
assign addr[39661]= -1844288924;
assign addr[39662]= -1803941934;
assign addr[39663]= -1761306505;
assign addr[39664]= -1716436725;
assign addr[39665]= -1669389513;
assign addr[39666]= -1620224553;
assign addr[39667]= -1569004214;
assign addr[39668]= -1515793473;
assign addr[39669]= -1460659832;
assign addr[39670]= -1403673233;
assign addr[39671]= -1344905966;
assign addr[39672]= -1284432584;
assign addr[39673]= -1222329801;
assign addr[39674]= -1158676398;
assign addr[39675]= -1093553126;
assign addr[39676]= -1027042599;
assign addr[39677]= -959229189;
assign addr[39678]= -890198924;
assign addr[39679]= -820039373;
assign addr[39680]= -748839539;
assign addr[39681]= -676689746;
assign addr[39682]= -603681519;
assign addr[39683]= -529907477;
assign addr[39684]= -455461206;
assign addr[39685]= -380437148;
assign addr[39686]= -304930476;
assign addr[39687]= -229036977;
assign addr[39688]= -152852926;
assign addr[39689]= -76474970;
assign addr[39690]= 0;
assign addr[39691]= 76474970;
assign addr[39692]= 152852926;
assign addr[39693]= 229036977;
assign addr[39694]= 304930476;
assign addr[39695]= 380437148;
assign addr[39696]= 455461206;
assign addr[39697]= 529907477;
assign addr[39698]= 603681519;
assign addr[39699]= 676689746;
assign addr[39700]= 748839539;
assign addr[39701]= 820039373;
assign addr[39702]= 890198924;
assign addr[39703]= 959229189;
assign addr[39704]= 1027042599;
assign addr[39705]= 1093553126;
assign addr[39706]= 1158676398;
assign addr[39707]= 1222329801;
assign addr[39708]= 1284432584;
assign addr[39709]= 1344905966;
assign addr[39710]= 1403673233;
assign addr[39711]= 1460659832;
assign addr[39712]= 1515793473;
assign addr[39713]= 1569004214;
assign addr[39714]= 1620224553;
assign addr[39715]= 1669389513;
assign addr[39716]= 1716436725;
assign addr[39717]= 1761306505;
assign addr[39718]= 1803941934;
assign addr[39719]= 1844288924;
assign addr[39720]= 1882296293;
assign addr[39721]= 1917915825;
assign addr[39722]= 1951102334;
assign addr[39723]= 1981813720;
assign addr[39724]= 2010011024;
assign addr[39725]= 2035658475;
assign addr[39726]= 2058723538;
assign addr[39727]= 2079176953;
assign addr[39728]= 2096992772;
assign addr[39729]= 2112148396;
assign addr[39730]= 2124624598;
assign addr[39731]= 2134405552;
assign addr[39732]= 2141478848;
assign addr[39733]= 2145835515;
assign addr[39734]= 2147470025;
assign addr[39735]= 2146380306;
assign addr[39736]= 2142567738;
assign addr[39737]= 2136037160;
assign addr[39738]= 2126796855;
assign addr[39739]= 2114858546;
assign addr[39740]= 2100237377;
assign addr[39741]= 2082951896;
assign addr[39742]= 2063024031;
assign addr[39743]= 2040479063;
assign addr[39744]= 2015345591;
assign addr[39745]= 1987655498;
assign addr[39746]= 1957443913;
assign addr[39747]= 1924749160;
assign addr[39748]= 1889612716;
assign addr[39749]= 1852079154;
assign addr[39750]= 1812196087;
assign addr[39751]= 1770014111;
assign addr[39752]= 1725586737;
assign addr[39753]= 1678970324;
assign addr[39754]= 1630224009;
assign addr[39755]= 1579409630;
assign addr[39756]= 1526591649;
assign addr[39757]= 1471837070;
assign addr[39758]= 1415215352;
assign addr[39759]= 1356798326;
assign addr[39760]= 1296660098;
assign addr[39761]= 1234876957;
assign addr[39762]= 1171527280;
assign addr[39763]= 1106691431;
assign addr[39764]= 1040451659;
assign addr[39765]= 972891995;
assign addr[39766]= 904098143;
assign addr[39767]= 834157373;
assign addr[39768]= 763158411;
assign addr[39769]= 691191324;
assign addr[39770]= 618347408;
assign addr[39771]= 544719071;
assign addr[39772]= 470399716;
assign addr[39773]= 395483624;
assign addr[39774]= 320065829;
assign addr[39775]= 244242007;
assign addr[39776]= 168108346;
assign addr[39777]= 91761426;
assign addr[39778]= 15298099;
assign addr[39779]= -61184634;
assign addr[39780]= -137589750;
assign addr[39781]= -213820322;
assign addr[39782]= -289779648;
assign addr[39783]= -365371365;
assign addr[39784]= -440499581;
assign addr[39785]= -515068990;
assign addr[39786]= -588984994;
assign addr[39787]= -662153826;
assign addr[39788]= -734482665;
assign addr[39789]= -805879757;
assign addr[39790]= -876254528;
assign addr[39791]= -945517704;
assign addr[39792]= -1013581418;
assign addr[39793]= -1080359326;
assign addr[39794]= -1145766716;
assign addr[39795]= -1209720613;
assign addr[39796]= -1272139887;
assign addr[39797]= -1332945355;
assign addr[39798]= -1392059879;
assign addr[39799]= -1449408469;
assign addr[39800]= -1504918373;
assign addr[39801]= -1558519173;
assign addr[39802]= -1610142873;
assign addr[39803]= -1659723983;
assign addr[39804]= -1707199606;
assign addr[39805]= -1752509516;
assign addr[39806]= -1795596234;
assign addr[39807]= -1836405100;
assign addr[39808]= -1874884346;
assign addr[39809]= -1910985158;
assign addr[39810]= -1944661739;
assign addr[39811]= -1975871368;
assign addr[39812]= -2004574453;
assign addr[39813]= -2030734582;
assign addr[39814]= -2054318569;
assign addr[39815]= -2075296495;
assign addr[39816]= -2093641749;
assign addr[39817]= -2109331059;
assign addr[39818]= -2122344521;
assign addr[39819]= -2132665626;
assign addr[39820]= -2140281282;
assign addr[39821]= -2145181827;
assign addr[39822]= -2147361045;
assign addr[39823]= -2146816171;
assign addr[39824]= -2143547897;
assign addr[39825]= -2137560369;
assign addr[39826]= -2128861181;
assign addr[39827]= -2117461370;
assign addr[39828]= -2103375398;
assign addr[39829]= -2086621133;
assign addr[39830]= -2067219829;
assign addr[39831]= -2045196100;
assign addr[39832]= -2020577882;
assign addr[39833]= -1993396407;
assign addr[39834]= -1963686155;
assign addr[39835]= -1931484818;
assign addr[39836]= -1896833245;
assign addr[39837]= -1859775393;
assign addr[39838]= -1820358275;
assign addr[39839]= -1778631892;
assign addr[39840]= -1734649179;
assign addr[39841]= -1688465931;
assign addr[39842]= -1640140734;
assign addr[39843]= -1589734894;
assign addr[39844]= -1537312353;
assign addr[39845]= -1482939614;
assign addr[39846]= -1426685652;
assign addr[39847]= -1368621831;
assign addr[39848]= -1308821808;
assign addr[39849]= -1247361445;
assign addr[39850]= -1184318708;
assign addr[39851]= -1119773573;
assign addr[39852]= -1053807919;
assign addr[39853]= -986505429;
assign addr[39854]= -917951481;
assign addr[39855]= -848233042;
assign addr[39856]= -777438554;
assign addr[39857]= -705657826;
assign addr[39858]= -632981917;
assign addr[39859]= -559503022;
assign addr[39860]= -485314355;
assign addr[39861]= -410510029;
assign addr[39862]= -335184940;
assign addr[39863]= -259434643;
assign addr[39864]= -183355234;
assign addr[39865]= -107043224;
assign addr[39866]= -30595422;
assign addr[39867]= 45891193;
assign addr[39868]= 122319591;
assign addr[39869]= 198592817;
assign addr[39870]= 274614114;
assign addr[39871]= 350287041;
assign addr[39872]= 425515602;
assign addr[39873]= 500204365;
assign addr[39874]= 574258580;
assign addr[39875]= 647584304;
assign addr[39876]= 720088517;
assign addr[39877]= 791679244;
assign addr[39878]= 862265664;
assign addr[39879]= 931758235;
assign addr[39880]= 1000068799;
assign addr[39881]= 1067110699;
assign addr[39882]= 1132798888;
assign addr[39883]= 1197050035;
assign addr[39884]= 1259782632;
assign addr[39885]= 1320917099;
assign addr[39886]= 1380375881;
assign addr[39887]= 1438083551;
assign addr[39888]= 1493966902;
assign addr[39889]= 1547955041;
assign addr[39890]= 1599979481;
assign addr[39891]= 1649974225;
assign addr[39892]= 1697875851;
assign addr[39893]= 1743623590;
assign addr[39894]= 1787159411;
assign addr[39895]= 1828428082;
assign addr[39896]= 1867377253;
assign addr[39897]= 1903957513;
assign addr[39898]= 1938122457;
assign addr[39899]= 1969828744;
assign addr[39900]= 1999036154;
assign addr[39901]= 2025707632;
assign addr[39902]= 2049809346;
assign addr[39903]= 2071310720;
assign addr[39904]= 2090184478;
assign addr[39905]= 2106406677;
assign addr[39906]= 2119956737;
assign addr[39907]= 2130817471;
assign addr[39908]= 2138975100;
assign addr[39909]= 2144419275;
assign addr[39910]= 2147143090;
assign addr[39911]= 2147143090;
assign addr[39912]= 2144419275;
assign addr[39913]= 2138975100;
assign addr[39914]= 2130817471;
assign addr[39915]= 2119956737;
assign addr[39916]= 2106406677;
assign addr[39917]= 2090184478;
assign addr[39918]= 2071310720;
assign addr[39919]= 2049809346;
assign addr[39920]= 2025707632;
assign addr[39921]= 1999036154;
assign addr[39922]= 1969828744;
assign addr[39923]= 1938122457;
assign addr[39924]= 1903957513;
assign addr[39925]= 1867377253;
assign addr[39926]= 1828428082;
assign addr[39927]= 1787159411;
assign addr[39928]= 1743623590;
assign addr[39929]= 1697875851;
assign addr[39930]= 1649974225;
assign addr[39931]= 1599979481;
assign addr[39932]= 1547955041;
assign addr[39933]= 1493966902;
assign addr[39934]= 1438083551;
assign addr[39935]= 1380375881;
assign addr[39936]= 1320917099;
assign addr[39937]= 1259782632;
assign addr[39938]= 1197050035;
assign addr[39939]= 1132798888;
assign addr[39940]= 1067110699;
assign addr[39941]= 1000068799;
assign addr[39942]= 931758235;
assign addr[39943]= 862265664;
assign addr[39944]= 791679244;
assign addr[39945]= 720088517;
assign addr[39946]= 647584304;
assign addr[39947]= 574258580;
assign addr[39948]= 500204365;
assign addr[39949]= 425515602;
assign addr[39950]= 350287041;
assign addr[39951]= 274614114;
assign addr[39952]= 198592817;
assign addr[39953]= 122319591;
assign addr[39954]= 45891193;
assign addr[39955]= -30595422;
assign addr[39956]= -107043224;
assign addr[39957]= -183355234;
assign addr[39958]= -259434643;
assign addr[39959]= -335184940;
assign addr[39960]= -410510029;
assign addr[39961]= -485314355;
assign addr[39962]= -559503022;
assign addr[39963]= -632981917;
assign addr[39964]= -705657826;
assign addr[39965]= -777438554;
assign addr[39966]= -848233042;
assign addr[39967]= -917951481;
assign addr[39968]= -986505429;
assign addr[39969]= -1053807919;
assign addr[39970]= -1119773573;
assign addr[39971]= -1184318708;
assign addr[39972]= -1247361445;
assign addr[39973]= -1308821808;
assign addr[39974]= -1368621831;
assign addr[39975]= -1426685652;
assign addr[39976]= -1482939614;
assign addr[39977]= -1537312353;
assign addr[39978]= -1589734894;
assign addr[39979]= -1640140734;
assign addr[39980]= -1688465931;
assign addr[39981]= -1734649179;
assign addr[39982]= -1778631892;
assign addr[39983]= -1820358275;
assign addr[39984]= -1859775393;
assign addr[39985]= -1896833245;
assign addr[39986]= -1931484818;
assign addr[39987]= -1963686155;
assign addr[39988]= -1993396407;
assign addr[39989]= -2020577882;
assign addr[39990]= -2045196100;
assign addr[39991]= -2067219829;
assign addr[39992]= -2086621133;
assign addr[39993]= -2103375398;
assign addr[39994]= -2117461370;
assign addr[39995]= -2128861181;
assign addr[39996]= -2137560369;
assign addr[39997]= -2143547897;
assign addr[39998]= -2146816171;
assign addr[39999]= -2147361045;
assign addr[40000]= -2145181827;
assign addr[40001]= -2140281282;
assign addr[40002]= -2132665626;
assign addr[40003]= -2122344521;
assign addr[40004]= -2109331059;
assign addr[40005]= -2093641749;
assign addr[40006]= -2075296495;
assign addr[40007]= -2054318569;
assign addr[40008]= -2030734582;
assign addr[40009]= -2004574453;
assign addr[40010]= -1975871368;
assign addr[40011]= -1944661739;
assign addr[40012]= -1910985158;
assign addr[40013]= -1874884346;
assign addr[40014]= -1836405100;
assign addr[40015]= -1795596234;
assign addr[40016]= -1752509516;
assign addr[40017]= -1707199606;
assign addr[40018]= -1659723983;
assign addr[40019]= -1610142873;
assign addr[40020]= -1558519173;
assign addr[40021]= -1504918373;
assign addr[40022]= -1449408469;
assign addr[40023]= -1392059879;
assign addr[40024]= -1332945355;
assign addr[40025]= -1272139887;
assign addr[40026]= -1209720613;
assign addr[40027]= -1145766716;
assign addr[40028]= -1080359326;
assign addr[40029]= -1013581418;
assign addr[40030]= -945517704;
assign addr[40031]= -876254528;
assign addr[40032]= -805879757;
assign addr[40033]= -734482665;
assign addr[40034]= -662153826;
assign addr[40035]= -588984994;
assign addr[40036]= -515068990;
assign addr[40037]= -440499581;
assign addr[40038]= -365371365;
assign addr[40039]= -289779648;
assign addr[40040]= -213820322;
assign addr[40041]= -137589750;
assign addr[40042]= -61184634;
assign addr[40043]= 15298099;
assign addr[40044]= 91761426;
assign addr[40045]= 168108346;
assign addr[40046]= 244242007;
assign addr[40047]= 320065829;
assign addr[40048]= 395483624;
assign addr[40049]= 470399716;
assign addr[40050]= 544719071;
assign addr[40051]= 618347408;
assign addr[40052]= 691191324;
assign addr[40053]= 763158411;
assign addr[40054]= 834157373;
assign addr[40055]= 904098143;
assign addr[40056]= 972891995;
assign addr[40057]= 1040451659;
assign addr[40058]= 1106691431;
assign addr[40059]= 1171527280;
assign addr[40060]= 1234876957;
assign addr[40061]= 1296660098;
assign addr[40062]= 1356798326;
assign addr[40063]= 1415215352;
assign addr[40064]= 1471837070;
assign addr[40065]= 1526591649;
assign addr[40066]= 1579409630;
assign addr[40067]= 1630224009;
assign addr[40068]= 1678970324;
assign addr[40069]= 1725586737;
assign addr[40070]= 1770014111;
assign addr[40071]= 1812196087;
assign addr[40072]= 1852079154;
assign addr[40073]= 1889612716;
assign addr[40074]= 1924749160;
assign addr[40075]= 1957443913;
assign addr[40076]= 1987655498;
assign addr[40077]= 2015345591;
assign addr[40078]= 2040479063;
assign addr[40079]= 2063024031;
assign addr[40080]= 2082951896;
assign addr[40081]= 2100237377;
assign addr[40082]= 2114858546;
assign addr[40083]= 2126796855;
assign addr[40084]= 2136037160;
assign addr[40085]= 2142567738;
assign addr[40086]= 2146380306;
assign addr[40087]= 2147470025;
assign addr[40088]= 2145835515;
assign addr[40089]= 2141478848;
assign addr[40090]= 2134405552;
assign addr[40091]= 2124624598;
assign addr[40092]= 2112148396;
assign addr[40093]= 2096992772;
assign addr[40094]= 2079176953;
assign addr[40095]= 2058723538;
assign addr[40096]= 2035658475;
assign addr[40097]= 2010011024;
assign addr[40098]= 1981813720;
assign addr[40099]= 1951102334;
assign addr[40100]= 1917915825;
assign addr[40101]= 1882296293;
assign addr[40102]= 1844288924;
assign addr[40103]= 1803941934;
assign addr[40104]= 1761306505;
assign addr[40105]= 1716436725;
assign addr[40106]= 1669389513;
assign addr[40107]= 1620224553;
assign addr[40108]= 1569004214;
assign addr[40109]= 1515793473;
assign addr[40110]= 1460659832;
assign addr[40111]= 1403673233;
assign addr[40112]= 1344905966;
assign addr[40113]= 1284432584;
assign addr[40114]= 1222329801;
assign addr[40115]= 1158676398;
assign addr[40116]= 1093553126;
assign addr[40117]= 1027042599;
assign addr[40118]= 959229189;
assign addr[40119]= 890198924;
assign addr[40120]= 820039373;
assign addr[40121]= 748839539;
assign addr[40122]= 676689746;
assign addr[40123]= 603681519;
assign addr[40124]= 529907477;
assign addr[40125]= 455461206;
assign addr[40126]= 380437148;
assign addr[40127]= 304930476;
assign addr[40128]= 229036977;
assign addr[40129]= 152852926;
assign addr[40130]= 76474970;
assign addr[40131]= 0;
assign addr[40132]= -76474970;
assign addr[40133]= -152852926;
assign addr[40134]= -229036977;
assign addr[40135]= -304930476;
assign addr[40136]= -380437148;
assign addr[40137]= -455461206;
assign addr[40138]= -529907477;
assign addr[40139]= -603681519;
assign addr[40140]= -676689746;
assign addr[40141]= -748839539;
assign addr[40142]= -820039373;
assign addr[40143]= -890198924;
assign addr[40144]= -959229189;
assign addr[40145]= -1027042599;
assign addr[40146]= -1093553126;
assign addr[40147]= -1158676398;
assign addr[40148]= -1222329801;
assign addr[40149]= -1284432584;
assign addr[40150]= -1344905966;
assign addr[40151]= -1403673233;
assign addr[40152]= -1460659832;
assign addr[40153]= -1515793473;
assign addr[40154]= -1569004214;
assign addr[40155]= -1620224553;
assign addr[40156]= -1669389513;
assign addr[40157]= -1716436725;
assign addr[40158]= -1761306505;
assign addr[40159]= -1803941934;
assign addr[40160]= -1844288924;
assign addr[40161]= -1882296293;
assign addr[40162]= -1917915825;
assign addr[40163]= -1951102334;
assign addr[40164]= -1981813720;
assign addr[40165]= -2010011024;
assign addr[40166]= -2035658475;
assign addr[40167]= -2058723538;
assign addr[40168]= -2079176953;
assign addr[40169]= -2096992772;
assign addr[40170]= -2112148396;
assign addr[40171]= -2124624598;
assign addr[40172]= -2134405552;
assign addr[40173]= -2141478848;
assign addr[40174]= -2145835515;
assign addr[40175]= -2147470025;
assign addr[40176]= -2146380306;
assign addr[40177]= -2142567738;
assign addr[40178]= -2136037160;
assign addr[40179]= -2126796855;
assign addr[40180]= -2114858546;
assign addr[40181]= -2100237377;
assign addr[40182]= -2082951896;
assign addr[40183]= -2063024031;
assign addr[40184]= -2040479063;
assign addr[40185]= -2015345591;
assign addr[40186]= -1987655498;
assign addr[40187]= -1957443913;
assign addr[40188]= -1924749160;
assign addr[40189]= -1889612716;
assign addr[40190]= -1852079154;
assign addr[40191]= -1812196087;
assign addr[40192]= -1770014111;
assign addr[40193]= -1725586737;
assign addr[40194]= -1678970324;
assign addr[40195]= -1630224009;
assign addr[40196]= -1579409630;
assign addr[40197]= -1526591649;
assign addr[40198]= -1471837070;
assign addr[40199]= -1415215352;
assign addr[40200]= -1356798326;
assign addr[40201]= -1296660098;
assign addr[40202]= -1234876957;
assign addr[40203]= -1171527280;
assign addr[40204]= -1106691431;
assign addr[40205]= -1040451659;
assign addr[40206]= -972891995;
assign addr[40207]= -904098143;
assign addr[40208]= -834157373;
assign addr[40209]= -763158411;
assign addr[40210]= -691191324;
assign addr[40211]= -618347408;
assign addr[40212]= -544719071;
assign addr[40213]= -470399716;
assign addr[40214]= -395483624;
assign addr[40215]= -320065829;
assign addr[40216]= -244242007;
assign addr[40217]= -168108346;
assign addr[40218]= -91761426;
assign addr[40219]= -15298099;
assign addr[40220]= 61184634;
assign addr[40221]= 137589750;
assign addr[40222]= 213820322;
assign addr[40223]= 289779648;
assign addr[40224]= 365371365;
assign addr[40225]= 440499581;
assign addr[40226]= 515068990;
assign addr[40227]= 588984994;
assign addr[40228]= 662153826;
assign addr[40229]= 734482665;
assign addr[40230]= 805879757;
assign addr[40231]= 876254528;
assign addr[40232]= 945517704;
assign addr[40233]= 1013581418;
assign addr[40234]= 1080359326;
assign addr[40235]= 1145766716;
assign addr[40236]= 1209720613;
assign addr[40237]= 1272139887;
assign addr[40238]= 1332945355;
assign addr[40239]= 1392059879;
assign addr[40240]= 1449408469;
assign addr[40241]= 1504918373;
assign addr[40242]= 1558519173;
assign addr[40243]= 1610142873;
assign addr[40244]= 1659723983;
assign addr[40245]= 1707199606;
assign addr[40246]= 1752509516;
assign addr[40247]= 1795596234;
assign addr[40248]= 1836405100;
assign addr[40249]= 1874884346;
assign addr[40250]= 1910985158;
assign addr[40251]= 1944661739;
assign addr[40252]= 1975871368;
assign addr[40253]= 2004574453;
assign addr[40254]= 2030734582;
assign addr[40255]= 2054318569;
assign addr[40256]= 2075296495;
assign addr[40257]= 2093641749;
assign addr[40258]= 2109331059;
assign addr[40259]= 2122344521;
assign addr[40260]= 2132665626;
assign addr[40261]= 2140281282;
assign addr[40262]= 2145181827;
assign addr[40263]= 2147361045;
assign addr[40264]= 2146816171;
assign addr[40265]= 2143547897;
assign addr[40266]= 2137560369;
assign addr[40267]= 2128861181;
assign addr[40268]= 2117461370;
assign addr[40269]= 2103375398;
assign addr[40270]= 2086621133;
assign addr[40271]= 2067219829;
assign addr[40272]= 2045196100;
assign addr[40273]= 2020577882;
assign addr[40274]= 1993396407;
assign addr[40275]= 1963686155;
assign addr[40276]= 1931484818;
assign addr[40277]= 1896833245;
assign addr[40278]= 1859775393;
assign addr[40279]= 1820358275;
assign addr[40280]= 1778631892;
assign addr[40281]= 1734649179;
assign addr[40282]= 1688465931;
assign addr[40283]= 1640140734;
assign addr[40284]= 1589734894;
assign addr[40285]= 1537312353;
assign addr[40286]= 1482939614;
assign addr[40287]= 1426685652;
assign addr[40288]= 1368621831;
assign addr[40289]= 1308821808;
assign addr[40290]= 1247361445;
assign addr[40291]= 1184318708;
assign addr[40292]= 1119773573;
assign addr[40293]= 1053807919;
assign addr[40294]= 986505429;
assign addr[40295]= 917951481;
assign addr[40296]= 848233042;
assign addr[40297]= 777438554;
assign addr[40298]= 705657826;
assign addr[40299]= 632981917;
assign addr[40300]= 559503022;
assign addr[40301]= 485314355;
assign addr[40302]= 410510029;
assign addr[40303]= 335184940;
assign addr[40304]= 259434643;
assign addr[40305]= 183355234;
assign addr[40306]= 107043224;
assign addr[40307]= 30595422;
assign addr[40308]= -45891193;
assign addr[40309]= -122319591;
assign addr[40310]= -198592817;
assign addr[40311]= -274614114;
assign addr[40312]= -350287041;
assign addr[40313]= -425515602;
assign addr[40314]= -500204365;
assign addr[40315]= -574258580;
assign addr[40316]= -647584304;
assign addr[40317]= -720088517;
assign addr[40318]= -791679244;
assign addr[40319]= -862265664;
assign addr[40320]= -931758235;
assign addr[40321]= -1000068799;
assign addr[40322]= -1067110699;
assign addr[40323]= -1132798888;
assign addr[40324]= -1197050035;
assign addr[40325]= -1259782632;
assign addr[40326]= -1320917099;
assign addr[40327]= -1380375881;
assign addr[40328]= -1438083551;
assign addr[40329]= -1493966902;
assign addr[40330]= -1547955041;
assign addr[40331]= -1599979481;
assign addr[40332]= -1649974225;
assign addr[40333]= -1697875851;
assign addr[40334]= -1743623590;
assign addr[40335]= -1787159411;
assign addr[40336]= -1828428082;
assign addr[40337]= -1867377253;
assign addr[40338]= -1903957513;
assign addr[40339]= -1938122457;
assign addr[40340]= -1969828744;
assign addr[40341]= -1999036154;
assign addr[40342]= -2025707632;
assign addr[40343]= -2049809346;
assign addr[40344]= -2071310720;
assign addr[40345]= -2090184478;
assign addr[40346]= -2106406677;
assign addr[40347]= -2119956737;
assign addr[40348]= -2130817471;
assign addr[40349]= -2138975100;
assign addr[40350]= -2144419275;
assign addr[40351]= -2147143090;
assign addr[40352]= -2147143090;
assign addr[40353]= -2144419275;
assign addr[40354]= -2138975100;
assign addr[40355]= -2130817471;
assign addr[40356]= -2119956737;
assign addr[40357]= -2106406677;
assign addr[40358]= -2090184478;
assign addr[40359]= -2071310720;
assign addr[40360]= -2049809346;
assign addr[40361]= -2025707632;
assign addr[40362]= -1999036154;
assign addr[40363]= -1969828744;
assign addr[40364]= -1938122457;
assign addr[40365]= -1903957513;
assign addr[40366]= -1867377253;
assign addr[40367]= -1828428082;
assign addr[40368]= -1787159411;
assign addr[40369]= -1743623590;
assign addr[40370]= -1697875851;
assign addr[40371]= -1649974225;
assign addr[40372]= -1599979481;
assign addr[40373]= -1547955041;
assign addr[40374]= -1493966902;
assign addr[40375]= -1438083551;
assign addr[40376]= -1380375881;
assign addr[40377]= -1320917099;
assign addr[40378]= -1259782632;
assign addr[40379]= -1197050035;
assign addr[40380]= -1132798888;
assign addr[40381]= -1067110699;
assign addr[40382]= -1000068799;
assign addr[40383]= -931758235;
assign addr[40384]= -862265664;
assign addr[40385]= -791679244;
assign addr[40386]= -720088517;
assign addr[40387]= -647584304;
assign addr[40388]= -574258580;
assign addr[40389]= -500204365;
assign addr[40390]= -425515602;
assign addr[40391]= -350287041;
assign addr[40392]= -274614114;
assign addr[40393]= -198592817;
assign addr[40394]= -122319591;
assign addr[40395]= -45891193;
assign addr[40396]= 30595422;
assign addr[40397]= 107043224;
assign addr[40398]= 183355234;
assign addr[40399]= 259434643;
assign addr[40400]= 335184940;
assign addr[40401]= 410510029;
assign addr[40402]= 485314355;
assign addr[40403]= 559503022;
assign addr[40404]= 632981917;
assign addr[40405]= 705657826;
assign addr[40406]= 777438554;
assign addr[40407]= 848233042;
assign addr[40408]= 917951481;
assign addr[40409]= 986505429;
assign addr[40410]= 1053807919;
assign addr[40411]= 1119773573;
assign addr[40412]= 1184318708;
assign addr[40413]= 1247361445;
assign addr[40414]= 1308821808;
assign addr[40415]= 1368621831;
assign addr[40416]= 1426685652;
assign addr[40417]= 1482939614;
assign addr[40418]= 1537312353;
assign addr[40419]= 1589734894;
assign addr[40420]= 1640140734;
assign addr[40421]= 1688465931;
assign addr[40422]= 1734649179;
assign addr[40423]= 1778631892;
assign addr[40424]= 1820358275;
assign addr[40425]= 1859775393;
assign addr[40426]= 1896833245;
assign addr[40427]= 1931484818;
assign addr[40428]= 1963686155;
assign addr[40429]= 1993396407;
assign addr[40430]= 2020577882;
assign addr[40431]= 2045196100;
assign addr[40432]= 2067219829;
assign addr[40433]= 2086621133;
assign addr[40434]= 2103375398;
assign addr[40435]= 2117461370;
assign addr[40436]= 2128861181;
assign addr[40437]= 2137560369;
assign addr[40438]= 2143547897;
assign addr[40439]= 2146816171;
assign addr[40440]= 2147361045;
assign addr[40441]= 2145181827;
assign addr[40442]= 2140281282;
assign addr[40443]= 2132665626;
assign addr[40444]= 2122344521;
assign addr[40445]= 2109331059;
assign addr[40446]= 2093641749;
assign addr[40447]= 2075296495;
assign addr[40448]= 2054318569;
assign addr[40449]= 2030734582;
assign addr[40450]= 2004574453;
assign addr[40451]= 1975871368;
assign addr[40452]= 1944661739;
assign addr[40453]= 1910985158;
assign addr[40454]= 1874884346;
assign addr[40455]= 1836405100;
assign addr[40456]= 1795596234;
assign addr[40457]= 1752509516;
assign addr[40458]= 1707199606;
assign addr[40459]= 1659723983;
assign addr[40460]= 1610142873;
assign addr[40461]= 1558519173;
assign addr[40462]= 1504918373;
assign addr[40463]= 1449408469;
assign addr[40464]= 1392059879;
assign addr[40465]= 1332945355;
assign addr[40466]= 1272139887;
assign addr[40467]= 1209720613;
assign addr[40468]= 1145766716;
assign addr[40469]= 1080359326;
assign addr[40470]= 1013581418;
assign addr[40471]= 945517704;
assign addr[40472]= 876254528;
assign addr[40473]= 805879757;
assign addr[40474]= 734482665;
assign addr[40475]= 662153826;
assign addr[40476]= 588984994;
assign addr[40477]= 515068990;
assign addr[40478]= 440499581;
assign addr[40479]= 365371365;
assign addr[40480]= 289779648;
assign addr[40481]= 213820322;
assign addr[40482]= 137589750;
assign addr[40483]= 61184634;
assign addr[40484]= -15298099;
assign addr[40485]= -91761426;
assign addr[40486]= -168108346;
assign addr[40487]= -244242007;
assign addr[40488]= -320065829;
assign addr[40489]= -395483624;
assign addr[40490]= -470399716;
assign addr[40491]= -544719071;
assign addr[40492]= -618347408;
assign addr[40493]= -691191324;
assign addr[40494]= -763158411;
assign addr[40495]= -834157373;
assign addr[40496]= -904098143;
assign addr[40497]= -972891995;
assign addr[40498]= -1040451659;
assign addr[40499]= -1106691431;
assign addr[40500]= -1171527280;
assign addr[40501]= -1234876957;
assign addr[40502]= -1296660098;
assign addr[40503]= -1356798326;
assign addr[40504]= -1415215352;
assign addr[40505]= -1471837070;
assign addr[40506]= -1526591649;
assign addr[40507]= -1579409630;
assign addr[40508]= -1630224009;
assign addr[40509]= -1678970324;
assign addr[40510]= -1725586737;
assign addr[40511]= -1770014111;
assign addr[40512]= -1812196087;
assign addr[40513]= -1852079154;
assign addr[40514]= -1889612716;
assign addr[40515]= -1924749160;
assign addr[40516]= -1957443913;
assign addr[40517]= -1987655498;
assign addr[40518]= -2015345591;
assign addr[40519]= -2040479063;
assign addr[40520]= -2063024031;
assign addr[40521]= -2082951896;
assign addr[40522]= -2100237377;
assign addr[40523]= -2114858546;
assign addr[40524]= -2126796855;
assign addr[40525]= -2136037160;
assign addr[40526]= -2142567738;
assign addr[40527]= -2146380306;
assign addr[40528]= -2147470025;
assign addr[40529]= -2145835515;
assign addr[40530]= -2141478848;
assign addr[40531]= -2134405552;
assign addr[40532]= -2124624598;
assign addr[40533]= -2112148396;
assign addr[40534]= -2096992772;
assign addr[40535]= -2079176953;
assign addr[40536]= -2058723538;
assign addr[40537]= -2035658475;
assign addr[40538]= -2010011024;
assign addr[40539]= -1981813720;
assign addr[40540]= -1951102334;
assign addr[40541]= -1917915825;
assign addr[40542]= -1882296293;
assign addr[40543]= -1844288924;
assign addr[40544]= -1803941934;
assign addr[40545]= -1761306505;
assign addr[40546]= -1716436725;
assign addr[40547]= -1669389513;
assign addr[40548]= -1620224553;
assign addr[40549]= -1569004214;
assign addr[40550]= -1515793473;
assign addr[40551]= -1460659832;
assign addr[40552]= -1403673233;
assign addr[40553]= -1344905966;
assign addr[40554]= -1284432584;
assign addr[40555]= -1222329801;
assign addr[40556]= -1158676398;
assign addr[40557]= -1093553126;
assign addr[40558]= -1027042599;
assign addr[40559]= -959229189;
assign addr[40560]= -890198924;
assign addr[40561]= -820039373;
assign addr[40562]= -748839539;
assign addr[40563]= -676689746;
assign addr[40564]= -603681519;
assign addr[40565]= -529907477;
assign addr[40566]= -455461206;
assign addr[40567]= -380437148;
assign addr[40568]= -304930476;
assign addr[40569]= -229036977;
assign addr[40570]= -152852926;
assign addr[40571]= -76474970;
assign addr[40572]= 0;
assign addr[40573]= 76474970;
assign addr[40574]= 152852926;
assign addr[40575]= 229036977;
assign addr[40576]= 304930476;
assign addr[40577]= 380437148;
assign addr[40578]= 455461206;
assign addr[40579]= 529907477;
assign addr[40580]= 603681519;
assign addr[40581]= 676689746;
assign addr[40582]= 748839539;
assign addr[40583]= 820039373;
assign addr[40584]= 890198924;
assign addr[40585]= 959229189;
assign addr[40586]= 1027042599;
assign addr[40587]= 1093553126;
assign addr[40588]= 1158676398;
assign addr[40589]= 1222329801;
assign addr[40590]= 1284432584;
assign addr[40591]= 1344905966;
assign addr[40592]= 1403673233;
assign addr[40593]= 1460659832;
assign addr[40594]= 1515793473;
assign addr[40595]= 1569004214;
assign addr[40596]= 1620224553;
assign addr[40597]= 1669389513;
assign addr[40598]= 1716436725;
assign addr[40599]= 1761306505;
assign addr[40600]= 1803941934;
assign addr[40601]= 1844288924;
assign addr[40602]= 1882296293;
assign addr[40603]= 1917915825;
assign addr[40604]= 1951102334;
assign addr[40605]= 1981813720;
assign addr[40606]= 2010011024;
assign addr[40607]= 2035658475;
assign addr[40608]= 2058723538;
assign addr[40609]= 2079176953;
assign addr[40610]= 2096992772;
assign addr[40611]= 2112148396;
assign addr[40612]= 2124624598;
assign addr[40613]= 2134405552;
assign addr[40614]= 2141478848;
assign addr[40615]= 2145835515;
assign addr[40616]= 2147470025;
assign addr[40617]= 2146380306;
assign addr[40618]= 2142567738;
assign addr[40619]= 2136037160;
assign addr[40620]= 2126796855;
assign addr[40621]= 2114858546;
assign addr[40622]= 2100237377;
assign addr[40623]= 2082951896;
assign addr[40624]= 2063024031;
assign addr[40625]= 2040479063;
assign addr[40626]= 2015345591;
assign addr[40627]= 1987655498;
assign addr[40628]= 1957443913;
assign addr[40629]= 1924749160;
assign addr[40630]= 1889612716;
assign addr[40631]= 1852079154;
assign addr[40632]= 1812196087;
assign addr[40633]= 1770014111;
assign addr[40634]= 1725586737;
assign addr[40635]= 1678970324;
assign addr[40636]= 1630224009;
assign addr[40637]= 1579409630;
assign addr[40638]= 1526591649;
assign addr[40639]= 1471837070;
assign addr[40640]= 1415215352;
assign addr[40641]= 1356798326;
assign addr[40642]= 1296660098;
assign addr[40643]= 1234876957;
assign addr[40644]= 1171527280;
assign addr[40645]= 1106691431;
assign addr[40646]= 1040451659;
assign addr[40647]= 972891995;
assign addr[40648]= 904098143;
assign addr[40649]= 834157373;
assign addr[40650]= 763158411;
assign addr[40651]= 691191324;
assign addr[40652]= 618347408;
assign addr[40653]= 544719071;
assign addr[40654]= 470399716;
assign addr[40655]= 395483624;
assign addr[40656]= 320065829;
assign addr[40657]= 244242007;
assign addr[40658]= 168108346;
assign addr[40659]= 91761426;
assign addr[40660]= 15298099;
assign addr[40661]= -61184634;
assign addr[40662]= -137589750;
assign addr[40663]= -213820322;
assign addr[40664]= -289779648;
assign addr[40665]= -365371365;
assign addr[40666]= -440499581;
assign addr[40667]= -515068990;
assign addr[40668]= -588984994;
assign addr[40669]= -662153826;
assign addr[40670]= -734482665;
assign addr[40671]= -805879757;
assign addr[40672]= -876254528;
assign addr[40673]= -945517704;
assign addr[40674]= -1013581418;
assign addr[40675]= -1080359326;
assign addr[40676]= -1145766716;
assign addr[40677]= -1209720613;
assign addr[40678]= -1272139887;
assign addr[40679]= -1332945355;
assign addr[40680]= -1392059879;
assign addr[40681]= -1449408469;
assign addr[40682]= -1504918373;
assign addr[40683]= -1558519173;
assign addr[40684]= -1610142873;
assign addr[40685]= -1659723983;
assign addr[40686]= -1707199606;
assign addr[40687]= -1752509516;
assign addr[40688]= -1795596234;
assign addr[40689]= -1836405100;
assign addr[40690]= -1874884346;
assign addr[40691]= -1910985158;
assign addr[40692]= -1944661739;
assign addr[40693]= -1975871368;
assign addr[40694]= -2004574453;
assign addr[40695]= -2030734582;
assign addr[40696]= -2054318569;
assign addr[40697]= -2075296495;
assign addr[40698]= -2093641749;
assign addr[40699]= -2109331059;
assign addr[40700]= -2122344521;
assign addr[40701]= -2132665626;
assign addr[40702]= -2140281282;
assign addr[40703]= -2145181827;
assign addr[40704]= -2147361045;
assign addr[40705]= -2146816171;
assign addr[40706]= -2143547897;
assign addr[40707]= -2137560369;
assign addr[40708]= -2128861181;
assign addr[40709]= -2117461370;
assign addr[40710]= -2103375398;
assign addr[40711]= -2086621133;
assign addr[40712]= -2067219829;
assign addr[40713]= -2045196100;
assign addr[40714]= -2020577882;
assign addr[40715]= -1993396407;
assign addr[40716]= -1963686155;
assign addr[40717]= -1931484818;
assign addr[40718]= -1896833245;
assign addr[40719]= -1859775393;
assign addr[40720]= -1820358275;
assign addr[40721]= -1778631892;
assign addr[40722]= -1734649179;
assign addr[40723]= -1688465931;
assign addr[40724]= -1640140734;
assign addr[40725]= -1589734894;
assign addr[40726]= -1537312353;
assign addr[40727]= -1482939614;
assign addr[40728]= -1426685652;
assign addr[40729]= -1368621831;
assign addr[40730]= -1308821808;
assign addr[40731]= -1247361445;
assign addr[40732]= -1184318708;
assign addr[40733]= -1119773573;
assign addr[40734]= -1053807919;
assign addr[40735]= -986505429;
assign addr[40736]= -917951481;
assign addr[40737]= -848233042;
assign addr[40738]= -777438554;
assign addr[40739]= -705657826;
assign addr[40740]= -632981917;
assign addr[40741]= -559503022;
assign addr[40742]= -485314355;
assign addr[40743]= -410510029;
assign addr[40744]= -335184940;
assign addr[40745]= -259434643;
assign addr[40746]= -183355234;
assign addr[40747]= -107043224;
assign addr[40748]= -30595422;
assign addr[40749]= 45891193;
assign addr[40750]= 122319591;
assign addr[40751]= 198592817;
assign addr[40752]= 274614114;
assign addr[40753]= 350287041;
assign addr[40754]= 425515602;
assign addr[40755]= 500204365;
assign addr[40756]= 574258580;
assign addr[40757]= 647584304;
assign addr[40758]= 720088517;
assign addr[40759]= 791679244;
assign addr[40760]= 862265664;
assign addr[40761]= 931758235;
assign addr[40762]= 1000068799;
assign addr[40763]= 1067110699;
assign addr[40764]= 1132798888;
assign addr[40765]= 1197050035;
assign addr[40766]= 1259782632;
assign addr[40767]= 1320917099;
assign addr[40768]= 1380375881;
assign addr[40769]= 1438083551;
assign addr[40770]= 1493966902;
assign addr[40771]= 1547955041;
assign addr[40772]= 1599979481;
assign addr[40773]= 1649974225;
assign addr[40774]= 1697875851;
assign addr[40775]= 1743623590;
assign addr[40776]= 1787159411;
assign addr[40777]= 1828428082;
assign addr[40778]= 1867377253;
assign addr[40779]= 1903957513;
assign addr[40780]= 1938122457;
assign addr[40781]= 1969828744;
assign addr[40782]= 1999036154;
assign addr[40783]= 2025707632;
assign addr[40784]= 2049809346;
assign addr[40785]= 2071310720;
assign addr[40786]= 2090184478;
assign addr[40787]= 2106406677;
assign addr[40788]= 2119956737;
assign addr[40789]= 2130817471;
assign addr[40790]= 2138975100;
assign addr[40791]= 2144419275;
assign addr[40792]= 2147143090;
assign addr[40793]= 2147143090;
assign addr[40794]= 2144419275;
assign addr[40795]= 2138975100;
assign addr[40796]= 2130817471;
assign addr[40797]= 2119956737;
assign addr[40798]= 2106406677;
assign addr[40799]= 2090184478;
assign addr[40800]= 2071310720;
assign addr[40801]= 2049809346;
assign addr[40802]= 2025707632;
assign addr[40803]= 1999036154;
assign addr[40804]= 1969828744;
assign addr[40805]= 1938122457;
assign addr[40806]= 1903957513;
assign addr[40807]= 1867377253;
assign addr[40808]= 1828428082;
assign addr[40809]= 1787159411;
assign addr[40810]= 1743623590;
assign addr[40811]= 1697875851;
assign addr[40812]= 1649974225;
assign addr[40813]= 1599979481;
assign addr[40814]= 1547955041;
assign addr[40815]= 1493966902;
assign addr[40816]= 1438083551;
assign addr[40817]= 1380375881;
assign addr[40818]= 1320917099;
assign addr[40819]= 1259782632;
assign addr[40820]= 1197050035;
assign addr[40821]= 1132798888;
assign addr[40822]= 1067110699;
assign addr[40823]= 1000068799;
assign addr[40824]= 931758235;
assign addr[40825]= 862265664;
assign addr[40826]= 791679244;
assign addr[40827]= 720088517;
assign addr[40828]= 647584304;
assign addr[40829]= 574258580;
assign addr[40830]= 500204365;
assign addr[40831]= 425515602;
assign addr[40832]= 350287041;
assign addr[40833]= 274614114;
assign addr[40834]= 198592817;
assign addr[40835]= 122319591;
assign addr[40836]= 45891193;
assign addr[40837]= -30595422;
assign addr[40838]= -107043224;
assign addr[40839]= -183355234;
assign addr[40840]= -259434643;
assign addr[40841]= -335184940;
assign addr[40842]= -410510029;
assign addr[40843]= -485314355;
assign addr[40844]= -559503022;
assign addr[40845]= -632981917;
assign addr[40846]= -705657826;
assign addr[40847]= -777438554;
assign addr[40848]= -848233042;
assign addr[40849]= -917951481;
assign addr[40850]= -986505429;
assign addr[40851]= -1053807919;
assign addr[40852]= -1119773573;
assign addr[40853]= -1184318708;
assign addr[40854]= -1247361445;
assign addr[40855]= -1308821808;
assign addr[40856]= -1368621831;
assign addr[40857]= -1426685652;
assign addr[40858]= -1482939614;
assign addr[40859]= -1537312353;
assign addr[40860]= -1589734894;
assign addr[40861]= -1640140734;
assign addr[40862]= -1688465931;
assign addr[40863]= -1734649179;
assign addr[40864]= -1778631892;
assign addr[40865]= -1820358275;
assign addr[40866]= -1859775393;
assign addr[40867]= -1896833245;
assign addr[40868]= -1931484818;
assign addr[40869]= -1963686155;
assign addr[40870]= -1993396407;
assign addr[40871]= -2020577882;
assign addr[40872]= -2045196100;
assign addr[40873]= -2067219829;
assign addr[40874]= -2086621133;
assign addr[40875]= -2103375398;
assign addr[40876]= -2117461370;
assign addr[40877]= -2128861181;
assign addr[40878]= -2137560369;
assign addr[40879]= -2143547897;
assign addr[40880]= -2146816171;
assign addr[40881]= -2147361045;
assign addr[40882]= -2145181827;
assign addr[40883]= -2140281282;
assign addr[40884]= -2132665626;
assign addr[40885]= -2122344521;
assign addr[40886]= -2109331059;
assign addr[40887]= -2093641749;
assign addr[40888]= -2075296495;
assign addr[40889]= -2054318569;
assign addr[40890]= -2030734582;
assign addr[40891]= -2004574453;
assign addr[40892]= -1975871368;
assign addr[40893]= -1944661739;
assign addr[40894]= -1910985158;
assign addr[40895]= -1874884346;
assign addr[40896]= -1836405100;
assign addr[40897]= -1795596234;
assign addr[40898]= -1752509516;
assign addr[40899]= -1707199606;
assign addr[40900]= -1659723983;
assign addr[40901]= -1610142873;
assign addr[40902]= -1558519173;
assign addr[40903]= -1504918373;
assign addr[40904]= -1449408469;
assign addr[40905]= -1392059879;
assign addr[40906]= -1332945355;
assign addr[40907]= -1272139887;
assign addr[40908]= -1209720613;
assign addr[40909]= -1145766716;
assign addr[40910]= -1080359326;
assign addr[40911]= -1013581418;
assign addr[40912]= -945517704;
assign addr[40913]= -876254528;
assign addr[40914]= -805879757;
assign addr[40915]= -734482665;
assign addr[40916]= -662153826;
assign addr[40917]= -588984994;
assign addr[40918]= -515068990;
assign addr[40919]= -440499581;
assign addr[40920]= -365371365;
assign addr[40921]= -289779648;
assign addr[40922]= -213820322;
assign addr[40923]= -137589750;
assign addr[40924]= -61184634;
assign addr[40925]= 15298099;
assign addr[40926]= 91761426;
assign addr[40927]= 168108346;
assign addr[40928]= 244242007;
assign addr[40929]= 320065829;
assign addr[40930]= 395483624;
assign addr[40931]= 470399716;
assign addr[40932]= 544719071;
assign addr[40933]= 618347408;
assign addr[40934]= 691191324;
assign addr[40935]= 763158411;
assign addr[40936]= 834157373;
assign addr[40937]= 904098143;
assign addr[40938]= 972891995;
assign addr[40939]= 1040451659;
assign addr[40940]= 1106691431;
assign addr[40941]= 1171527280;
assign addr[40942]= 1234876957;
assign addr[40943]= 1296660098;
assign addr[40944]= 1356798326;
assign addr[40945]= 1415215352;
assign addr[40946]= 1471837070;
assign addr[40947]= 1526591649;
assign addr[40948]= 1579409630;
assign addr[40949]= 1630224009;
assign addr[40950]= 1678970324;
assign addr[40951]= 1725586737;
assign addr[40952]= 1770014111;
assign addr[40953]= 1812196087;
assign addr[40954]= 1852079154;
assign addr[40955]= 1889612716;
assign addr[40956]= 1924749160;
assign addr[40957]= 1957443913;
assign addr[40958]= 1987655498;
assign addr[40959]= 2015345591;
assign addr[40960]= 2040479063;
assign addr[40961]= 2063024031;
assign addr[40962]= 2082951896;
assign addr[40963]= 2100237377;
assign addr[40964]= 2114858546;
assign addr[40965]= 2126796855;
assign addr[40966]= 2136037160;
assign addr[40967]= 2142567738;
assign addr[40968]= 2146380306;
assign addr[40969]= 2147470025;
assign addr[40970]= 2145835515;
assign addr[40971]= 2141478848;
assign addr[40972]= 2134405552;
assign addr[40973]= 2124624598;
assign addr[40974]= 2112148396;
assign addr[40975]= 2096992772;
assign addr[40976]= 2079176953;
assign addr[40977]= 2058723538;
assign addr[40978]= 2035658475;
assign addr[40979]= 2010011024;
assign addr[40980]= 1981813720;
assign addr[40981]= 1951102334;
assign addr[40982]= 1917915825;
assign addr[40983]= 1882296293;
assign addr[40984]= 1844288924;
assign addr[40985]= 1803941934;
assign addr[40986]= 1761306505;
assign addr[40987]= 1716436725;
assign addr[40988]= 1669389513;
assign addr[40989]= 1620224553;
assign addr[40990]= 1569004214;
assign addr[40991]= 1515793473;
assign addr[40992]= 1460659832;
assign addr[40993]= 1403673233;
assign addr[40994]= 1344905966;
assign addr[40995]= 1284432584;
assign addr[40996]= 1222329801;
assign addr[40997]= 1158676398;
assign addr[40998]= 1093553126;
assign addr[40999]= 1027042599;
assign addr[41000]= 959229189;
assign addr[41001]= 890198924;
assign addr[41002]= 820039373;
assign addr[41003]= 748839539;
assign addr[41004]= 676689746;
assign addr[41005]= 603681519;
assign addr[41006]= 529907477;
assign addr[41007]= 455461206;
assign addr[41008]= 380437148;
assign addr[41009]= 304930476;
assign addr[41010]= 229036977;
assign addr[41011]= 152852926;
assign addr[41012]= 76474970;
assign addr[41013]= 0;
assign addr[41014]= -76474970;
assign addr[41015]= -152852926;
assign addr[41016]= -229036977;
assign addr[41017]= -304930476;
assign addr[41018]= -380437148;
assign addr[41019]= -455461206;
assign addr[41020]= -529907477;
assign addr[41021]= -603681519;
assign addr[41022]= -676689746;
assign addr[41023]= -748839539;
assign addr[41024]= -820039373;
assign addr[41025]= -890198924;
assign addr[41026]= -959229189;
assign addr[41027]= -1027042599;
assign addr[41028]= -1093553126;
assign addr[41029]= -1158676398;
assign addr[41030]= -1222329801;
assign addr[41031]= -1284432584;
assign addr[41032]= -1344905966;
assign addr[41033]= -1403673233;
assign addr[41034]= -1460659832;
assign addr[41035]= -1515793473;
assign addr[41036]= -1569004214;
assign addr[41037]= -1620224553;
assign addr[41038]= -1669389513;
assign addr[41039]= -1716436725;
assign addr[41040]= -1761306505;
assign addr[41041]= -1803941934;
assign addr[41042]= -1844288924;
assign addr[41043]= -1882296293;
assign addr[41044]= -1917915825;
assign addr[41045]= -1951102334;
assign addr[41046]= -1981813720;
assign addr[41047]= -2010011024;
assign addr[41048]= -2035658475;
assign addr[41049]= -2058723538;
assign addr[41050]= -2079176953;
assign addr[41051]= -2096992772;
assign addr[41052]= -2112148396;
assign addr[41053]= -2124624598;
assign addr[41054]= -2134405552;
assign addr[41055]= -2141478848;
assign addr[41056]= -2145835515;
assign addr[41057]= -2147470025;
assign addr[41058]= -2146380306;
assign addr[41059]= -2142567738;
assign addr[41060]= -2136037160;
assign addr[41061]= -2126796855;
assign addr[41062]= -2114858546;
assign addr[41063]= -2100237377;
assign addr[41064]= -2082951896;
assign addr[41065]= -2063024031;
assign addr[41066]= -2040479063;
assign addr[41067]= -2015345591;
assign addr[41068]= -1987655498;
assign addr[41069]= -1957443913;
assign addr[41070]= -1924749160;
assign addr[41071]= -1889612716;
assign addr[41072]= -1852079154;
assign addr[41073]= -1812196087;
assign addr[41074]= -1770014111;
assign addr[41075]= -1725586737;
assign addr[41076]= -1678970324;
assign addr[41077]= -1630224009;
assign addr[41078]= -1579409630;
assign addr[41079]= -1526591649;
assign addr[41080]= -1471837070;
assign addr[41081]= -1415215352;
assign addr[41082]= -1356798326;
assign addr[41083]= -1296660098;
assign addr[41084]= -1234876957;
assign addr[41085]= -1171527280;
assign addr[41086]= -1106691431;
assign addr[41087]= -1040451659;
assign addr[41088]= -972891995;
assign addr[41089]= -904098143;
assign addr[41090]= -834157373;
assign addr[41091]= -763158411;
assign addr[41092]= -691191324;
assign addr[41093]= -618347408;
assign addr[41094]= -544719071;
assign addr[41095]= -470399716;
assign addr[41096]= -395483624;
assign addr[41097]= -320065829;
assign addr[41098]= -244242007;
assign addr[41099]= -168108346;
assign addr[41100]= -91761426;
assign addr[41101]= -15298099;
assign addr[41102]= 61184634;
assign addr[41103]= 137589750;
assign addr[41104]= 213820322;
assign addr[41105]= 289779648;
assign addr[41106]= 365371365;
assign addr[41107]= 440499581;
assign addr[41108]= 515068990;
assign addr[41109]= 588984994;
assign addr[41110]= 662153826;
assign addr[41111]= 734482665;
assign addr[41112]= 805879757;
assign addr[41113]= 876254528;
assign addr[41114]= 945517704;
assign addr[41115]= 1013581418;
assign addr[41116]= 1080359326;
assign addr[41117]= 1145766716;
assign addr[41118]= 1209720613;
assign addr[41119]= 1272139887;
assign addr[41120]= 1332945355;
assign addr[41121]= 1392059879;
assign addr[41122]= 1449408469;
assign addr[41123]= 1504918373;
assign addr[41124]= 1558519173;
assign addr[41125]= 1610142873;
assign addr[41126]= 1659723983;
assign addr[41127]= 1707199606;
assign addr[41128]= 1752509516;
assign addr[41129]= 1795596234;
assign addr[41130]= 1836405100;
assign addr[41131]= 1874884346;
assign addr[41132]= 1910985158;
assign addr[41133]= 1944661739;
assign addr[41134]= 1975871368;
assign addr[41135]= 2004574453;
assign addr[41136]= 2030734582;
assign addr[41137]= 2054318569;
assign addr[41138]= 2075296495;
assign addr[41139]= 2093641749;
assign addr[41140]= 2109331059;
assign addr[41141]= 2122344521;
assign addr[41142]= 2132665626;
assign addr[41143]= 2140281282;
assign addr[41144]= 2145181827;
assign addr[41145]= 2147361045;
assign addr[41146]= 2146816171;
assign addr[41147]= 2143547897;
assign addr[41148]= 2137560369;
assign addr[41149]= 2128861181;
assign addr[41150]= 2117461370;
assign addr[41151]= 2103375398;
assign addr[41152]= 2086621133;
assign addr[41153]= 2067219829;
assign addr[41154]= 2045196100;
assign addr[41155]= 2020577882;
assign addr[41156]= 1993396407;
assign addr[41157]= 1963686155;
assign addr[41158]= 1931484818;
assign addr[41159]= 1896833245;
assign addr[41160]= 1859775393;
assign addr[41161]= 1820358275;
assign addr[41162]= 1778631892;
assign addr[41163]= 1734649179;
assign addr[41164]= 1688465931;
assign addr[41165]= 1640140734;
assign addr[41166]= 1589734894;
assign addr[41167]= 1537312353;
assign addr[41168]= 1482939614;
assign addr[41169]= 1426685652;
assign addr[41170]= 1368621831;
assign addr[41171]= 1308821808;
assign addr[41172]= 1247361445;
assign addr[41173]= 1184318708;
assign addr[41174]= 1119773573;
assign addr[41175]= 1053807919;
assign addr[41176]= 986505429;
assign addr[41177]= 917951481;
assign addr[41178]= 848233042;
assign addr[41179]= 777438554;
assign addr[41180]= 705657826;
assign addr[41181]= 632981917;
assign addr[41182]= 559503022;
assign addr[41183]= 485314355;
assign addr[41184]= 410510029;
assign addr[41185]= 335184940;
assign addr[41186]= 259434643;
assign addr[41187]= 183355234;
assign addr[41188]= 107043224;
assign addr[41189]= 30595422;
assign addr[41190]= -45891193;
assign addr[41191]= -122319591;
assign addr[41192]= -198592817;
assign addr[41193]= -274614114;
assign addr[41194]= -350287041;
assign addr[41195]= -425515602;
assign addr[41196]= -500204365;
assign addr[41197]= -574258580;
assign addr[41198]= -647584304;
assign addr[41199]= -720088517;
assign addr[41200]= -791679244;
assign addr[41201]= -862265664;
assign addr[41202]= -931758235;
assign addr[41203]= -1000068799;
assign addr[41204]= -1067110699;
assign addr[41205]= -1132798888;
assign addr[41206]= -1197050035;
assign addr[41207]= -1259782632;
assign addr[41208]= -1320917099;
assign addr[41209]= -1380375881;
assign addr[41210]= -1438083551;
assign addr[41211]= -1493966902;
assign addr[41212]= -1547955041;
assign addr[41213]= -1599979481;
assign addr[41214]= -1649974225;
assign addr[41215]= -1697875851;
assign addr[41216]= -1743623590;
assign addr[41217]= -1787159411;
assign addr[41218]= -1828428082;
assign addr[41219]= -1867377253;
assign addr[41220]= -1903957513;
assign addr[41221]= -1938122457;
assign addr[41222]= -1969828744;
assign addr[41223]= -1999036154;
assign addr[41224]= -2025707632;
assign addr[41225]= -2049809346;
assign addr[41226]= -2071310720;
assign addr[41227]= -2090184478;
assign addr[41228]= -2106406677;
assign addr[41229]= -2119956737;
assign addr[41230]= -2130817471;
assign addr[41231]= -2138975100;
assign addr[41232]= -2144419275;
assign addr[41233]= -2147143090;
assign addr[41234]= -2147143090;
assign addr[41235]= -2144419275;
assign addr[41236]= -2138975100;
assign addr[41237]= -2130817471;
assign addr[41238]= -2119956737;
assign addr[41239]= -2106406677;
assign addr[41240]= -2090184478;
assign addr[41241]= -2071310720;
assign addr[41242]= -2049809346;
assign addr[41243]= -2025707632;
assign addr[41244]= -1999036154;
assign addr[41245]= -1969828744;
assign addr[41246]= -1938122457;
assign addr[41247]= -1903957513;
assign addr[41248]= -1867377253;
assign addr[41249]= -1828428082;
assign addr[41250]= -1787159411;
assign addr[41251]= -1743623590;
assign addr[41252]= -1697875851;
assign addr[41253]= -1649974225;
assign addr[41254]= -1599979481;
assign addr[41255]= -1547955041;
assign addr[41256]= -1493966902;
assign addr[41257]= -1438083551;
assign addr[41258]= -1380375881;
assign addr[41259]= -1320917099;
assign addr[41260]= -1259782632;
assign addr[41261]= -1197050035;
assign addr[41262]= -1132798888;
assign addr[41263]= -1067110699;
assign addr[41264]= -1000068799;
assign addr[41265]= -931758235;
assign addr[41266]= -862265664;
assign addr[41267]= -791679244;
assign addr[41268]= -720088517;
assign addr[41269]= -647584304;
assign addr[41270]= -574258580;
assign addr[41271]= -500204365;
assign addr[41272]= -425515602;
assign addr[41273]= -350287041;
assign addr[41274]= -274614114;
assign addr[41275]= -198592817;
assign addr[41276]= -122319591;
assign addr[41277]= -45891193;
assign addr[41278]= 30595422;
assign addr[41279]= 107043224;
assign addr[41280]= 183355234;
assign addr[41281]= 259434643;
assign addr[41282]= 335184940;
assign addr[41283]= 410510029;
assign addr[41284]= 485314355;
assign addr[41285]= 559503022;
assign addr[41286]= 632981917;
assign addr[41287]= 705657826;
assign addr[41288]= 777438554;
assign addr[41289]= 848233042;
assign addr[41290]= 917951481;
assign addr[41291]= 986505429;
assign addr[41292]= 1053807919;
assign addr[41293]= 1119773573;
assign addr[41294]= 1184318708;
assign addr[41295]= 1247361445;
assign addr[41296]= 1308821808;
assign addr[41297]= 1368621831;
assign addr[41298]= 1426685652;
assign addr[41299]= 1482939614;
assign addr[41300]= 1537312353;
assign addr[41301]= 1589734894;
assign addr[41302]= 1640140734;
assign addr[41303]= 1688465931;
assign addr[41304]= 1734649179;
assign addr[41305]= 1778631892;
assign addr[41306]= 1820358275;
assign addr[41307]= 1859775393;
assign addr[41308]= 1896833245;
assign addr[41309]= 1931484818;
assign addr[41310]= 1963686155;
assign addr[41311]= 1993396407;
assign addr[41312]= 2020577882;
assign addr[41313]= 2045196100;
assign addr[41314]= 2067219829;
assign addr[41315]= 2086621133;
assign addr[41316]= 2103375398;
assign addr[41317]= 2117461370;
assign addr[41318]= 2128861181;
assign addr[41319]= 2137560369;
assign addr[41320]= 2143547897;
assign addr[41321]= 2146816171;
assign addr[41322]= 2147361045;
assign addr[41323]= 2145181827;
assign addr[41324]= 2140281282;
assign addr[41325]= 2132665626;
assign addr[41326]= 2122344521;
assign addr[41327]= 2109331059;
assign addr[41328]= 2093641749;
assign addr[41329]= 2075296495;
assign addr[41330]= 2054318569;
assign addr[41331]= 2030734582;
assign addr[41332]= 2004574453;
assign addr[41333]= 1975871368;
assign addr[41334]= 1944661739;
assign addr[41335]= 1910985158;
assign addr[41336]= 1874884346;
assign addr[41337]= 1836405100;
assign addr[41338]= 1795596234;
assign addr[41339]= 1752509516;
assign addr[41340]= 1707199606;
assign addr[41341]= 1659723983;
assign addr[41342]= 1610142873;
assign addr[41343]= 1558519173;
assign addr[41344]= 1504918373;
assign addr[41345]= 1449408469;
assign addr[41346]= 1392059879;
assign addr[41347]= 1332945355;
assign addr[41348]= 1272139887;
assign addr[41349]= 1209720613;
assign addr[41350]= 1145766716;
assign addr[41351]= 1080359326;
assign addr[41352]= 1013581418;
assign addr[41353]= 945517704;
assign addr[41354]= 876254528;
assign addr[41355]= 805879757;
assign addr[41356]= 734482665;
assign addr[41357]= 662153826;
assign addr[41358]= 588984994;
assign addr[41359]= 515068990;
assign addr[41360]= 440499581;
assign addr[41361]= 365371365;
assign addr[41362]= 289779648;
assign addr[41363]= 213820322;
assign addr[41364]= 137589750;
assign addr[41365]= 61184634;
assign addr[41366]= -15298099;
assign addr[41367]= -91761426;
assign addr[41368]= -168108346;
assign addr[41369]= -244242007;
assign addr[41370]= -320065829;
assign addr[41371]= -395483624;
assign addr[41372]= -470399716;
assign addr[41373]= -544719071;
assign addr[41374]= -618347408;
assign addr[41375]= -691191324;
assign addr[41376]= -763158411;
assign addr[41377]= -834157373;
assign addr[41378]= -904098143;
assign addr[41379]= -972891995;
assign addr[41380]= -1040451659;
assign addr[41381]= -1106691431;
assign addr[41382]= -1171527280;
assign addr[41383]= -1234876957;
assign addr[41384]= -1296660098;
assign addr[41385]= -1356798326;
assign addr[41386]= -1415215352;
assign addr[41387]= -1471837070;
assign addr[41388]= -1526591649;
assign addr[41389]= -1579409630;
assign addr[41390]= -1630224009;
assign addr[41391]= -1678970324;
assign addr[41392]= -1725586737;
assign addr[41393]= -1770014111;
assign addr[41394]= -1812196087;
assign addr[41395]= -1852079154;
assign addr[41396]= -1889612716;
assign addr[41397]= -1924749160;
assign addr[41398]= -1957443913;
assign addr[41399]= -1987655498;
assign addr[41400]= -2015345591;
assign addr[41401]= -2040479063;
assign addr[41402]= -2063024031;
assign addr[41403]= -2082951896;
assign addr[41404]= -2100237377;
assign addr[41405]= -2114858546;
assign addr[41406]= -2126796855;
assign addr[41407]= -2136037160;
assign addr[41408]= -2142567738;
assign addr[41409]= -2146380306;
assign addr[41410]= -2147470025;
assign addr[41411]= -2145835515;
assign addr[41412]= -2141478848;
assign addr[41413]= -2134405552;
assign addr[41414]= -2124624598;
assign addr[41415]= -2112148396;
assign addr[41416]= -2096992772;
assign addr[41417]= -2079176953;
assign addr[41418]= -2058723538;
assign addr[41419]= -2035658475;
assign addr[41420]= -2010011024;
assign addr[41421]= -1981813720;
assign addr[41422]= -1951102334;
assign addr[41423]= -1917915825;
assign addr[41424]= -1882296293;
assign addr[41425]= -1844288924;
assign addr[41426]= -1803941934;
assign addr[41427]= -1761306505;
assign addr[41428]= -1716436725;
assign addr[41429]= -1669389513;
assign addr[41430]= -1620224553;
assign addr[41431]= -1569004214;
assign addr[41432]= -1515793473;
assign addr[41433]= -1460659832;
assign addr[41434]= -1403673233;
assign addr[41435]= -1344905966;
assign addr[41436]= -1284432584;
assign addr[41437]= -1222329801;
assign addr[41438]= -1158676398;
assign addr[41439]= -1093553126;
assign addr[41440]= -1027042599;
assign addr[41441]= -959229189;
assign addr[41442]= -890198924;
assign addr[41443]= -820039373;
assign addr[41444]= -748839539;
assign addr[41445]= -676689746;
assign addr[41446]= -603681519;
assign addr[41447]= -529907477;
assign addr[41448]= -455461206;
assign addr[41449]= -380437148;
assign addr[41450]= -304930476;
assign addr[41451]= -229036977;
assign addr[41452]= -152852926;
assign addr[41453]= -76474970;
assign addr[41454]= 0;
assign addr[41455]= 76474970;
assign addr[41456]= 152852926;
assign addr[41457]= 229036977;
assign addr[41458]= 304930476;
assign addr[41459]= 380437148;
assign addr[41460]= 455461206;
assign addr[41461]= 529907477;
assign addr[41462]= 603681519;
assign addr[41463]= 676689746;
assign addr[41464]= 748839539;
assign addr[41465]= 820039373;
assign addr[41466]= 890198924;
assign addr[41467]= 959229189;
assign addr[41468]= 1027042599;
assign addr[41469]= 1093553126;
assign addr[41470]= 1158676398;
assign addr[41471]= 1222329801;
assign addr[41472]= 1284432584;
assign addr[41473]= 1344905966;
assign addr[41474]= 1403673233;
assign addr[41475]= 1460659832;
assign addr[41476]= 1515793473;
assign addr[41477]= 1569004214;
assign addr[41478]= 1620224553;
assign addr[41479]= 1669389513;
assign addr[41480]= 1716436725;
assign addr[41481]= 1761306505;
assign addr[41482]= 1803941934;
assign addr[41483]= 1844288924;
assign addr[41484]= 1882296293;
assign addr[41485]= 1917915825;
assign addr[41486]= 1951102334;
assign addr[41487]= 1981813720;
assign addr[41488]= 2010011024;
assign addr[41489]= 2035658475;
assign addr[41490]= 2058723538;
assign addr[41491]= 2079176953;
assign addr[41492]= 2096992772;
assign addr[41493]= 2112148396;
assign addr[41494]= 2124624598;
assign addr[41495]= 2134405552;
assign addr[41496]= 2141478848;
assign addr[41497]= 2145835515;
assign addr[41498]= 2147470025;
assign addr[41499]= 2146380306;
assign addr[41500]= 2142567738;
assign addr[41501]= 2136037160;
assign addr[41502]= 2126796855;
assign addr[41503]= 2114858546;
assign addr[41504]= 2100237377;
assign addr[41505]= 2082951896;
assign addr[41506]= 2063024031;
assign addr[41507]= 2040479063;
assign addr[41508]= 2015345591;
assign addr[41509]= 1987655498;
assign addr[41510]= 1957443913;
assign addr[41511]= 1924749160;
assign addr[41512]= 1889612716;
assign addr[41513]= 1852079154;
assign addr[41514]= 1812196087;
assign addr[41515]= 1770014111;
assign addr[41516]= 1725586737;
assign addr[41517]= 1678970324;
assign addr[41518]= 1630224009;
assign addr[41519]= 1579409630;
assign addr[41520]= 1526591649;
assign addr[41521]= 1471837070;
assign addr[41522]= 1415215352;
assign addr[41523]= 1356798326;
assign addr[41524]= 1296660098;
assign addr[41525]= 1234876957;
assign addr[41526]= 1171527280;
assign addr[41527]= 1106691431;
assign addr[41528]= 1040451659;
assign addr[41529]= 972891995;
assign addr[41530]= 904098143;
assign addr[41531]= 834157373;
assign addr[41532]= 763158411;
assign addr[41533]= 691191324;
assign addr[41534]= 618347408;
assign addr[41535]= 544719071;
assign addr[41536]= 470399716;
assign addr[41537]= 395483624;
assign addr[41538]= 320065829;
assign addr[41539]= 244242007;
assign addr[41540]= 168108346;
assign addr[41541]= 91761426;
assign addr[41542]= 15298099;
assign addr[41543]= -61184634;
assign addr[41544]= -137589750;
assign addr[41545]= -213820322;
assign addr[41546]= -289779648;
assign addr[41547]= -365371365;
assign addr[41548]= -440499581;
assign addr[41549]= -515068990;
assign addr[41550]= -588984994;
assign addr[41551]= -662153826;
assign addr[41552]= -734482665;
assign addr[41553]= -805879757;
assign addr[41554]= -876254528;
assign addr[41555]= -945517704;
assign addr[41556]= -1013581418;
assign addr[41557]= -1080359326;
assign addr[41558]= -1145766716;
assign addr[41559]= -1209720613;
assign addr[41560]= -1272139887;
assign addr[41561]= -1332945355;
assign addr[41562]= -1392059879;
assign addr[41563]= -1449408469;
assign addr[41564]= -1504918373;
assign addr[41565]= -1558519173;
assign addr[41566]= -1610142873;
assign addr[41567]= -1659723983;
assign addr[41568]= -1707199606;
assign addr[41569]= -1752509516;
assign addr[41570]= -1795596234;
assign addr[41571]= -1836405100;
assign addr[41572]= -1874884346;
assign addr[41573]= -1910985158;
assign addr[41574]= -1944661739;
assign addr[41575]= -1975871368;
assign addr[41576]= -2004574453;
assign addr[41577]= -2030734582;
assign addr[41578]= -2054318569;
assign addr[41579]= -2075296495;
assign addr[41580]= -2093641749;
assign addr[41581]= -2109331059;
assign addr[41582]= -2122344521;
assign addr[41583]= -2132665626;
assign addr[41584]= -2140281282;
assign addr[41585]= -2145181827;
assign addr[41586]= -2147361045;
assign addr[41587]= -2146816171;
assign addr[41588]= -2143547897;
assign addr[41589]= -2137560369;
assign addr[41590]= -2128861181;
assign addr[41591]= -2117461370;
assign addr[41592]= -2103375398;
assign addr[41593]= -2086621133;
assign addr[41594]= -2067219829;
assign addr[41595]= -2045196100;
assign addr[41596]= -2020577882;
assign addr[41597]= -1993396407;
assign addr[41598]= -1963686155;
assign addr[41599]= -1931484818;
assign addr[41600]= -1896833245;
assign addr[41601]= -1859775393;
assign addr[41602]= -1820358275;
assign addr[41603]= -1778631892;
assign addr[41604]= -1734649179;
assign addr[41605]= -1688465931;
assign addr[41606]= -1640140734;
assign addr[41607]= -1589734894;
assign addr[41608]= -1537312353;
assign addr[41609]= -1482939614;
assign addr[41610]= -1426685652;
assign addr[41611]= -1368621831;
assign addr[41612]= -1308821808;
assign addr[41613]= -1247361445;
assign addr[41614]= -1184318708;
assign addr[41615]= -1119773573;
assign addr[41616]= -1053807919;
assign addr[41617]= -986505429;
assign addr[41618]= -917951481;
assign addr[41619]= -848233042;
assign addr[41620]= -777438554;
assign addr[41621]= -705657826;
assign addr[41622]= -632981917;
assign addr[41623]= -559503022;
assign addr[41624]= -485314355;
assign addr[41625]= -410510029;
assign addr[41626]= -335184940;
assign addr[41627]= -259434643;
assign addr[41628]= -183355234;
assign addr[41629]= -107043224;
assign addr[41630]= -30595422;
assign addr[41631]= 45891193;
assign addr[41632]= 122319591;
assign addr[41633]= 198592817;
assign addr[41634]= 274614114;
assign addr[41635]= 350287041;
assign addr[41636]= 425515602;
assign addr[41637]= 500204365;
assign addr[41638]= 574258580;
assign addr[41639]= 647584304;
assign addr[41640]= 720088517;
assign addr[41641]= 791679244;
assign addr[41642]= 862265664;
assign addr[41643]= 931758235;
assign addr[41644]= 1000068799;
assign addr[41645]= 1067110699;
assign addr[41646]= 1132798888;
assign addr[41647]= 1197050035;
assign addr[41648]= 1259782632;
assign addr[41649]= 1320917099;
assign addr[41650]= 1380375881;
assign addr[41651]= 1438083551;
assign addr[41652]= 1493966902;
assign addr[41653]= 1547955041;
assign addr[41654]= 1599979481;
assign addr[41655]= 1649974225;
assign addr[41656]= 1697875851;
assign addr[41657]= 1743623590;
assign addr[41658]= 1787159411;
assign addr[41659]= 1828428082;
assign addr[41660]= 1867377253;
assign addr[41661]= 1903957513;
assign addr[41662]= 1938122457;
assign addr[41663]= 1969828744;
assign addr[41664]= 1999036154;
assign addr[41665]= 2025707632;
assign addr[41666]= 2049809346;
assign addr[41667]= 2071310720;
assign addr[41668]= 2090184478;
assign addr[41669]= 2106406677;
assign addr[41670]= 2119956737;
assign addr[41671]= 2130817471;
assign addr[41672]= 2138975100;
assign addr[41673]= 2144419275;
assign addr[41674]= 2147143090;
assign addr[41675]= 2147143090;
assign addr[41676]= 2144419275;
assign addr[41677]= 2138975100;
assign addr[41678]= 2130817471;
assign addr[41679]= 2119956737;
assign addr[41680]= 2106406677;
assign addr[41681]= 2090184478;
assign addr[41682]= 2071310720;
assign addr[41683]= 2049809346;
assign addr[41684]= 2025707632;
assign addr[41685]= 1999036154;
assign addr[41686]= 1969828744;
assign addr[41687]= 1938122457;
assign addr[41688]= 1903957513;
assign addr[41689]= 1867377253;
assign addr[41690]= 1828428082;
assign addr[41691]= 1787159411;
assign addr[41692]= 1743623590;
assign addr[41693]= 1697875851;
assign addr[41694]= 1649974225;
assign addr[41695]= 1599979481;
assign addr[41696]= 1547955041;
assign addr[41697]= 1493966902;
assign addr[41698]= 1438083551;
assign addr[41699]= 1380375881;
assign addr[41700]= 1320917099;
assign addr[41701]= 1259782632;
assign addr[41702]= 1197050035;
assign addr[41703]= 1132798888;
assign addr[41704]= 1067110699;
assign addr[41705]= 1000068799;
assign addr[41706]= 931758235;
assign addr[41707]= 862265664;
assign addr[41708]= 791679244;
assign addr[41709]= 720088517;
assign addr[41710]= 647584304;
assign addr[41711]= 574258580;
assign addr[41712]= 500204365;
assign addr[41713]= 425515602;
assign addr[41714]= 350287041;
assign addr[41715]= 274614114;
assign addr[41716]= 198592817;
assign addr[41717]= 122319591;
assign addr[41718]= 45891193;
assign addr[41719]= -30595422;
assign addr[41720]= -107043224;
assign addr[41721]= -183355234;
assign addr[41722]= -259434643;
assign addr[41723]= -335184940;
assign addr[41724]= -410510029;
assign addr[41725]= -485314355;
assign addr[41726]= -559503022;
assign addr[41727]= -632981917;
assign addr[41728]= -705657826;
assign addr[41729]= -777438554;
assign addr[41730]= -848233042;
assign addr[41731]= -917951481;
assign addr[41732]= -986505429;
assign addr[41733]= -1053807919;
assign addr[41734]= -1119773573;
assign addr[41735]= -1184318708;
assign addr[41736]= -1247361445;
assign addr[41737]= -1308821808;
assign addr[41738]= -1368621831;
assign addr[41739]= -1426685652;
assign addr[41740]= -1482939614;
assign addr[41741]= -1537312353;
assign addr[41742]= -1589734894;
assign addr[41743]= -1640140734;
assign addr[41744]= -1688465931;
assign addr[41745]= -1734649179;
assign addr[41746]= -1778631892;
assign addr[41747]= -1820358275;
assign addr[41748]= -1859775393;
assign addr[41749]= -1896833245;
assign addr[41750]= -1931484818;
assign addr[41751]= -1963686155;
assign addr[41752]= -1993396407;
assign addr[41753]= -2020577882;
assign addr[41754]= -2045196100;
assign addr[41755]= -2067219829;
assign addr[41756]= -2086621133;
assign addr[41757]= -2103375398;
assign addr[41758]= -2117461370;
assign addr[41759]= -2128861181;
assign addr[41760]= -2137560369;
assign addr[41761]= -2143547897;
assign addr[41762]= -2146816171;
assign addr[41763]= -2147361045;
assign addr[41764]= -2145181827;
assign addr[41765]= -2140281282;
assign addr[41766]= -2132665626;
assign addr[41767]= -2122344521;
assign addr[41768]= -2109331059;
assign addr[41769]= -2093641749;
assign addr[41770]= -2075296495;
assign addr[41771]= -2054318569;
assign addr[41772]= -2030734582;
assign addr[41773]= -2004574453;
assign addr[41774]= -1975871368;
assign addr[41775]= -1944661739;
assign addr[41776]= -1910985158;
assign addr[41777]= -1874884346;
assign addr[41778]= -1836405100;
assign addr[41779]= -1795596234;
assign addr[41780]= -1752509516;
assign addr[41781]= -1707199606;
assign addr[41782]= -1659723983;
assign addr[41783]= -1610142873;
assign addr[41784]= -1558519173;
assign addr[41785]= -1504918373;
assign addr[41786]= -1449408469;
assign addr[41787]= -1392059879;
assign addr[41788]= -1332945355;
assign addr[41789]= -1272139887;
assign addr[41790]= -1209720613;
assign addr[41791]= -1145766716;
assign addr[41792]= -1080359326;
assign addr[41793]= -1013581418;
assign addr[41794]= -945517704;
assign addr[41795]= -876254528;
assign addr[41796]= -805879757;
assign addr[41797]= -734482665;
assign addr[41798]= -662153826;
assign addr[41799]= -588984994;
assign addr[41800]= -515068990;
assign addr[41801]= -440499581;
assign addr[41802]= -365371365;
assign addr[41803]= -289779648;
assign addr[41804]= -213820322;
assign addr[41805]= -137589750;
assign addr[41806]= -61184634;
assign addr[41807]= 15298099;
assign addr[41808]= 91761426;
assign addr[41809]= 168108346;
assign addr[41810]= 244242007;
assign addr[41811]= 320065829;
assign addr[41812]= 395483624;
assign addr[41813]= 470399716;
assign addr[41814]= 544719071;
assign addr[41815]= 618347408;
assign addr[41816]= 691191324;
assign addr[41817]= 763158411;
assign addr[41818]= 834157373;
assign addr[41819]= 904098143;
assign addr[41820]= 972891995;
assign addr[41821]= 1040451659;
assign addr[41822]= 1106691431;
assign addr[41823]= 1171527280;
assign addr[41824]= 1234876957;
assign addr[41825]= 1296660098;
assign addr[41826]= 1356798326;
assign addr[41827]= 1415215352;
assign addr[41828]= 1471837070;
assign addr[41829]= 1526591649;
assign addr[41830]= 1579409630;
assign addr[41831]= 1630224009;
assign addr[41832]= 1678970324;
assign addr[41833]= 1725586737;
assign addr[41834]= 1770014111;
assign addr[41835]= 1812196087;
assign addr[41836]= 1852079154;
assign addr[41837]= 1889612716;
assign addr[41838]= 1924749160;
assign addr[41839]= 1957443913;
assign addr[41840]= 1987655498;
assign addr[41841]= 2015345591;
assign addr[41842]= 2040479063;
assign addr[41843]= 2063024031;
assign addr[41844]= 2082951896;
assign addr[41845]= 2100237377;
assign addr[41846]= 2114858546;
assign addr[41847]= 2126796855;
assign addr[41848]= 2136037160;
assign addr[41849]= 2142567738;
assign addr[41850]= 2146380306;
assign addr[41851]= 2147470025;
assign addr[41852]= 2145835515;
assign addr[41853]= 2141478848;
assign addr[41854]= 2134405552;
assign addr[41855]= 2124624598;
assign addr[41856]= 2112148396;
assign addr[41857]= 2096992772;
assign addr[41858]= 2079176953;
assign addr[41859]= 2058723538;
assign addr[41860]= 2035658475;
assign addr[41861]= 2010011024;
assign addr[41862]= 1981813720;
assign addr[41863]= 1951102334;
assign addr[41864]= 1917915825;
assign addr[41865]= 1882296293;
assign addr[41866]= 1844288924;
assign addr[41867]= 1803941934;
assign addr[41868]= 1761306505;
assign addr[41869]= 1716436725;
assign addr[41870]= 1669389513;
assign addr[41871]= 1620224553;
assign addr[41872]= 1569004214;
assign addr[41873]= 1515793473;
assign addr[41874]= 1460659832;
assign addr[41875]= 1403673233;
assign addr[41876]= 1344905966;
assign addr[41877]= 1284432584;
assign addr[41878]= 1222329801;
assign addr[41879]= 1158676398;
assign addr[41880]= 1093553126;
assign addr[41881]= 1027042599;
assign addr[41882]= 959229189;
assign addr[41883]= 890198924;
assign addr[41884]= 820039373;
assign addr[41885]= 748839539;
assign addr[41886]= 676689746;
assign addr[41887]= 603681519;
assign addr[41888]= 529907477;
assign addr[41889]= 455461206;
assign addr[41890]= 380437148;
assign addr[41891]= 304930476;
assign addr[41892]= 229036977;
assign addr[41893]= 152852926;
assign addr[41894]= 76474970;
assign addr[41895]= 0;
assign addr[41896]= -76474970;
assign addr[41897]= -152852926;
assign addr[41898]= -229036977;
assign addr[41899]= -304930476;
assign addr[41900]= -380437148;
assign addr[41901]= -455461206;
assign addr[41902]= -529907477;
assign addr[41903]= -603681519;
assign addr[41904]= -676689746;
assign addr[41905]= -748839539;
assign addr[41906]= -820039373;
assign addr[41907]= -890198924;
assign addr[41908]= -959229189;
assign addr[41909]= -1027042599;
assign addr[41910]= -1093553126;
assign addr[41911]= -1158676398;
assign addr[41912]= -1222329801;
assign addr[41913]= -1284432584;
assign addr[41914]= -1344905966;
assign addr[41915]= -1403673233;
assign addr[41916]= -1460659832;
assign addr[41917]= -1515793473;
assign addr[41918]= -1569004214;
assign addr[41919]= -1620224553;
assign addr[41920]= -1669389513;
assign addr[41921]= -1716436725;
assign addr[41922]= -1761306505;
assign addr[41923]= -1803941934;
assign addr[41924]= -1844288924;
assign addr[41925]= -1882296293;
assign addr[41926]= -1917915825;
assign addr[41927]= -1951102334;
assign addr[41928]= -1981813720;
assign addr[41929]= -2010011024;
assign addr[41930]= -2035658475;
assign addr[41931]= -2058723538;
assign addr[41932]= -2079176953;
assign addr[41933]= -2096992772;
assign addr[41934]= -2112148396;
assign addr[41935]= -2124624598;
assign addr[41936]= -2134405552;
assign addr[41937]= -2141478848;
assign addr[41938]= -2145835515;
assign addr[41939]= -2147470025;
assign addr[41940]= -2146380306;
assign addr[41941]= -2142567738;
assign addr[41942]= -2136037160;
assign addr[41943]= -2126796855;
assign addr[41944]= -2114858546;
assign addr[41945]= -2100237377;
assign addr[41946]= -2082951896;
assign addr[41947]= -2063024031;
assign addr[41948]= -2040479063;
assign addr[41949]= -2015345591;
assign addr[41950]= -1987655498;
assign addr[41951]= -1957443913;
assign addr[41952]= -1924749160;
assign addr[41953]= -1889612716;
assign addr[41954]= -1852079154;
assign addr[41955]= -1812196087;
assign addr[41956]= -1770014111;
assign addr[41957]= -1725586737;
assign addr[41958]= -1678970324;
assign addr[41959]= -1630224009;
assign addr[41960]= -1579409630;
assign addr[41961]= -1526591649;
assign addr[41962]= -1471837070;
assign addr[41963]= -1415215352;
assign addr[41964]= -1356798326;
assign addr[41965]= -1296660098;
assign addr[41966]= -1234876957;
assign addr[41967]= -1171527280;
assign addr[41968]= -1106691431;
assign addr[41969]= -1040451659;
assign addr[41970]= -972891995;
assign addr[41971]= -904098143;
assign addr[41972]= -834157373;
assign addr[41973]= -763158411;
assign addr[41974]= -691191324;
assign addr[41975]= -618347408;
assign addr[41976]= -544719071;
assign addr[41977]= -470399716;
assign addr[41978]= -395483624;
assign addr[41979]= -320065829;
assign addr[41980]= -244242007;
assign addr[41981]= -168108346;
assign addr[41982]= -91761426;
assign addr[41983]= -15298099;
assign addr[41984]= 61184634;
assign addr[41985]= 137589750;
assign addr[41986]= 213820322;
assign addr[41987]= 289779648;
assign addr[41988]= 365371365;
assign addr[41989]= 440499581;
assign addr[41990]= 515068990;
assign addr[41991]= 588984994;
assign addr[41992]= 662153826;
assign addr[41993]= 734482665;
assign addr[41994]= 805879757;
assign addr[41995]= 876254528;
assign addr[41996]= 945517704;
assign addr[41997]= 1013581418;
assign addr[41998]= 1080359326;
assign addr[41999]= 1145766716;
assign addr[42000]= 1209720613;
assign addr[42001]= 1272139887;
assign addr[42002]= 1332945355;
assign addr[42003]= 1392059879;
assign addr[42004]= 1449408469;
assign addr[42005]= 1504918373;
assign addr[42006]= 1558519173;
assign addr[42007]= 1610142873;
assign addr[42008]= 1659723983;
assign addr[42009]= 1707199606;
assign addr[42010]= 1752509516;
assign addr[42011]= 1795596234;
assign addr[42012]= 1836405100;
assign addr[42013]= 1874884346;
assign addr[42014]= 1910985158;
assign addr[42015]= 1944661739;
assign addr[42016]= 1975871368;
assign addr[42017]= 2004574453;
assign addr[42018]= 2030734582;
assign addr[42019]= 2054318569;
assign addr[42020]= 2075296495;
assign addr[42021]= 2093641749;
assign addr[42022]= 2109331059;
assign addr[42023]= 2122344521;
assign addr[42024]= 2132665626;
assign addr[42025]= 2140281282;
assign addr[42026]= 2145181827;
assign addr[42027]= 2147361045;
assign addr[42028]= 2146816171;
assign addr[42029]= 2143547897;
assign addr[42030]= 2137560369;
assign addr[42031]= 2128861181;
assign addr[42032]= 2117461370;
assign addr[42033]= 2103375398;
assign addr[42034]= 2086621133;
assign addr[42035]= 2067219829;
assign addr[42036]= 2045196100;
assign addr[42037]= 2020577882;
assign addr[42038]= 1993396407;
assign addr[42039]= 1963686155;
assign addr[42040]= 1931484818;
assign addr[42041]= 1896833245;
assign addr[42042]= 1859775393;
assign addr[42043]= 1820358275;
assign addr[42044]= 1778631892;
assign addr[42045]= 1734649179;
assign addr[42046]= 1688465931;
assign addr[42047]= 1640140734;
assign addr[42048]= 1589734894;
assign addr[42049]= 1537312353;
assign addr[42050]= 1482939614;
assign addr[42051]= 1426685652;
assign addr[42052]= 1368621831;
assign addr[42053]= 1308821808;
assign addr[42054]= 1247361445;
assign addr[42055]= 1184318708;
assign addr[42056]= 1119773573;
assign addr[42057]= 1053807919;
assign addr[42058]= 986505429;
assign addr[42059]= 917951481;
assign addr[42060]= 848233042;
assign addr[42061]= 777438554;
assign addr[42062]= 705657826;
assign addr[42063]= 632981917;
assign addr[42064]= 559503022;
assign addr[42065]= 485314355;
assign addr[42066]= 410510029;
assign addr[42067]= 335184940;
assign addr[42068]= 259434643;
assign addr[42069]= 183355234;
assign addr[42070]= 107043224;
assign addr[42071]= 30595422;
assign addr[42072]= -45891193;
assign addr[42073]= -122319591;
assign addr[42074]= -198592817;
assign addr[42075]= -274614114;
assign addr[42076]= -350287041;
assign addr[42077]= -425515602;
assign addr[42078]= -500204365;
assign addr[42079]= -574258580;
assign addr[42080]= -647584304;
assign addr[42081]= -720088517;
assign addr[42082]= -791679244;
assign addr[42083]= -862265664;
assign addr[42084]= -931758235;
assign addr[42085]= -1000068799;
assign addr[42086]= -1067110699;
assign addr[42087]= -1132798888;
assign addr[42088]= -1197050035;
assign addr[42089]= -1259782632;
assign addr[42090]= -1320917099;
assign addr[42091]= -1380375881;
assign addr[42092]= -1438083551;
assign addr[42093]= -1493966902;
assign addr[42094]= -1547955041;
assign addr[42095]= -1599979481;
assign addr[42096]= -1649974225;
assign addr[42097]= -1697875851;
assign addr[42098]= -1743623590;
assign addr[42099]= -1787159411;
assign addr[42100]= -1828428082;
assign addr[42101]= -1867377253;
assign addr[42102]= -1903957513;
assign addr[42103]= -1938122457;
assign addr[42104]= -1969828744;
assign addr[42105]= -1999036154;
assign addr[42106]= -2025707632;
assign addr[42107]= -2049809346;
assign addr[42108]= -2071310720;
assign addr[42109]= -2090184478;
assign addr[42110]= -2106406677;
assign addr[42111]= -2119956737;
assign addr[42112]= -2130817471;
assign addr[42113]= -2138975100;
assign addr[42114]= -2144419275;
assign addr[42115]= -2147143090;
assign addr[42116]= -2147143090;
assign addr[42117]= -2144419275;
assign addr[42118]= -2138975100;
assign addr[42119]= -2130817471;
assign addr[42120]= -2119956737;
assign addr[42121]= -2106406677;
assign addr[42122]= -2090184478;
assign addr[42123]= -2071310720;
assign addr[42124]= -2049809346;
assign addr[42125]= -2025707632;
assign addr[42126]= -1999036154;
assign addr[42127]= -1969828744;
assign addr[42128]= -1938122457;
assign addr[42129]= -1903957513;
assign addr[42130]= -1867377253;
assign addr[42131]= -1828428082;
assign addr[42132]= -1787159411;
assign addr[42133]= -1743623590;
assign addr[42134]= -1697875851;
assign addr[42135]= -1649974225;
assign addr[42136]= -1599979481;
assign addr[42137]= -1547955041;
assign addr[42138]= -1493966902;
assign addr[42139]= -1438083551;
assign addr[42140]= -1380375881;
assign addr[42141]= -1320917099;
assign addr[42142]= -1259782632;
assign addr[42143]= -1197050035;
assign addr[42144]= -1132798888;
assign addr[42145]= -1067110699;
assign addr[42146]= -1000068799;
assign addr[42147]= -931758235;
assign addr[42148]= -862265664;
assign addr[42149]= -791679244;
assign addr[42150]= -720088517;
assign addr[42151]= -647584304;
assign addr[42152]= -574258580;
assign addr[42153]= -500204365;
assign addr[42154]= -425515602;
assign addr[42155]= -350287041;
assign addr[42156]= -274614114;
assign addr[42157]= -198592817;
assign addr[42158]= -122319591;
assign addr[42159]= -45891193;
assign addr[42160]= 30595422;
assign addr[42161]= 107043224;
assign addr[42162]= 183355234;
assign addr[42163]= 259434643;
assign addr[42164]= 335184940;
assign addr[42165]= 410510029;
assign addr[42166]= 485314355;
assign addr[42167]= 559503022;
assign addr[42168]= 632981917;
assign addr[42169]= 705657826;
assign addr[42170]= 777438554;
assign addr[42171]= 848233042;
assign addr[42172]= 917951481;
assign addr[42173]= 986505429;
assign addr[42174]= 1053807919;
assign addr[42175]= 1119773573;
assign addr[42176]= 1184318708;
assign addr[42177]= 1247361445;
assign addr[42178]= 1308821808;
assign addr[42179]= 1368621831;
assign addr[42180]= 1426685652;
assign addr[42181]= 1482939614;
assign addr[42182]= 1537312353;
assign addr[42183]= 1589734894;
assign addr[42184]= 1640140734;
assign addr[42185]= 1688465931;
assign addr[42186]= 1734649179;
assign addr[42187]= 1778631892;
assign addr[42188]= 1820358275;
assign addr[42189]= 1859775393;
assign addr[42190]= 1896833245;
assign addr[42191]= 1931484818;
assign addr[42192]= 1963686155;
assign addr[42193]= 1993396407;
assign addr[42194]= 2020577882;
assign addr[42195]= 2045196100;
assign addr[42196]= 2067219829;
assign addr[42197]= 2086621133;
assign addr[42198]= 2103375398;
assign addr[42199]= 2117461370;
assign addr[42200]= 2128861181;
assign addr[42201]= 2137560369;
assign addr[42202]= 2143547897;
assign addr[42203]= 2146816171;
assign addr[42204]= 2147361045;
assign addr[42205]= 2145181827;
assign addr[42206]= 2140281282;
assign addr[42207]= 2132665626;
assign addr[42208]= 2122344521;
assign addr[42209]= 2109331059;
assign addr[42210]= 2093641749;
assign addr[42211]= 2075296495;
assign addr[42212]= 2054318569;
assign addr[42213]= 2030734582;
assign addr[42214]= 2004574453;
assign addr[42215]= 1975871368;
assign addr[42216]= 1944661739;
assign addr[42217]= 1910985158;
assign addr[42218]= 1874884346;
assign addr[42219]= 1836405100;
assign addr[42220]= 1795596234;
assign addr[42221]= 1752509516;
assign addr[42222]= 1707199606;
assign addr[42223]= 1659723983;
assign addr[42224]= 1610142873;
assign addr[42225]= 1558519173;
assign addr[42226]= 1504918373;
assign addr[42227]= 1449408469;
assign addr[42228]= 1392059879;
assign addr[42229]= 1332945355;
assign addr[42230]= 1272139887;
assign addr[42231]= 1209720613;
assign addr[42232]= 1145766716;
assign addr[42233]= 1080359326;
assign addr[42234]= 1013581418;
assign addr[42235]= 945517704;
assign addr[42236]= 876254528;
assign addr[42237]= 805879757;
assign addr[42238]= 734482665;
assign addr[42239]= 662153826;
assign addr[42240]= 588984994;
assign addr[42241]= 515068990;
assign addr[42242]= 440499581;
assign addr[42243]= 365371365;
assign addr[42244]= 289779648;
assign addr[42245]= 213820322;
assign addr[42246]= 137589750;
assign addr[42247]= 61184634;
assign addr[42248]= -15298099;
assign addr[42249]= -91761426;
assign addr[42250]= -168108346;
assign addr[42251]= -244242007;
assign addr[42252]= -320065829;
assign addr[42253]= -395483624;
assign addr[42254]= -470399716;
assign addr[42255]= -544719071;
assign addr[42256]= -618347408;
assign addr[42257]= -691191324;
assign addr[42258]= -763158411;
assign addr[42259]= -834157373;
assign addr[42260]= -904098143;
assign addr[42261]= -972891995;
assign addr[42262]= -1040451659;
assign addr[42263]= -1106691431;
assign addr[42264]= -1171527280;
assign addr[42265]= -1234876957;
assign addr[42266]= -1296660098;
assign addr[42267]= -1356798326;
assign addr[42268]= -1415215352;
assign addr[42269]= -1471837070;
assign addr[42270]= -1526591649;
assign addr[42271]= -1579409630;
assign addr[42272]= -1630224009;
assign addr[42273]= -1678970324;
assign addr[42274]= -1725586737;
assign addr[42275]= -1770014111;
assign addr[42276]= -1812196087;
assign addr[42277]= -1852079154;
assign addr[42278]= -1889612716;
assign addr[42279]= -1924749160;
assign addr[42280]= -1957443913;
assign addr[42281]= -1987655498;
assign addr[42282]= -2015345591;
assign addr[42283]= -2040479063;
assign addr[42284]= -2063024031;
assign addr[42285]= -2082951896;
assign addr[42286]= -2100237377;
assign addr[42287]= -2114858546;
assign addr[42288]= -2126796855;
assign addr[42289]= -2136037160;
assign addr[42290]= -2142567738;
assign addr[42291]= -2146380306;
assign addr[42292]= -2147470025;
assign addr[42293]= -2145835515;
assign addr[42294]= -2141478848;
assign addr[42295]= -2134405552;
assign addr[42296]= -2124624598;
assign addr[42297]= -2112148396;
assign addr[42298]= -2096992772;
assign addr[42299]= -2079176953;
assign addr[42300]= -2058723538;
assign addr[42301]= -2035658475;
assign addr[42302]= -2010011024;
assign addr[42303]= -1981813720;
assign addr[42304]= -1951102334;
assign addr[42305]= -1917915825;
assign addr[42306]= -1882296293;
assign addr[42307]= -1844288924;
assign addr[42308]= -1803941934;
assign addr[42309]= -1761306505;
assign addr[42310]= -1716436725;
assign addr[42311]= -1669389513;
assign addr[42312]= -1620224553;
assign addr[42313]= -1569004214;
assign addr[42314]= -1515793473;
assign addr[42315]= -1460659832;
assign addr[42316]= -1403673233;
assign addr[42317]= -1344905966;
assign addr[42318]= -1284432584;
assign addr[42319]= -1222329801;
assign addr[42320]= -1158676398;
assign addr[42321]= -1093553126;
assign addr[42322]= -1027042599;
assign addr[42323]= -959229189;
assign addr[42324]= -890198924;
assign addr[42325]= -820039373;
assign addr[42326]= -748839539;
assign addr[42327]= -676689746;
assign addr[42328]= -603681519;
assign addr[42329]= -529907477;
assign addr[42330]= -455461206;
assign addr[42331]= -380437148;
assign addr[42332]= -304930476;
assign addr[42333]= -229036977;
assign addr[42334]= -152852926;
assign addr[42335]= -76474970;
assign addr[42336]= 0;
assign addr[42337]= 76474970;
assign addr[42338]= 152852926;
assign addr[42339]= 229036977;
assign addr[42340]= 304930476;
assign addr[42341]= 380437148;
assign addr[42342]= 455461206;
assign addr[42343]= 529907477;
assign addr[42344]= 603681519;
assign addr[42345]= 676689746;
assign addr[42346]= 748839539;
assign addr[42347]= 820039373;
assign addr[42348]= 890198924;
assign addr[42349]= 959229189;
assign addr[42350]= 1027042599;
assign addr[42351]= 1093553126;
assign addr[42352]= 1158676398;
assign addr[42353]= 1222329801;
assign addr[42354]= 1284432584;
assign addr[42355]= 1344905966;
assign addr[42356]= 1403673233;
assign addr[42357]= 1460659832;
assign addr[42358]= 1515793473;
assign addr[42359]= 1569004214;
assign addr[42360]= 1620224553;
assign addr[42361]= 1669389513;
assign addr[42362]= 1716436725;
assign addr[42363]= 1761306505;
assign addr[42364]= 1803941934;
assign addr[42365]= 1844288924;
assign addr[42366]= 1882296293;
assign addr[42367]= 1917915825;
assign addr[42368]= 1951102334;
assign addr[42369]= 1981813720;
assign addr[42370]= 2010011024;
assign addr[42371]= 2035658475;
assign addr[42372]= 2058723538;
assign addr[42373]= 2079176953;
assign addr[42374]= 2096992772;
assign addr[42375]= 2112148396;
assign addr[42376]= 2124624598;
assign addr[42377]= 2134405552;
assign addr[42378]= 2141478848;
assign addr[42379]= 2145835515;
assign addr[42380]= 2147470025;
assign addr[42381]= 2146380306;
assign addr[42382]= 2142567738;
assign addr[42383]= 2136037160;
assign addr[42384]= 2126796855;
assign addr[42385]= 2114858546;
assign addr[42386]= 2100237377;
assign addr[42387]= 2082951896;
assign addr[42388]= 2063024031;
assign addr[42389]= 2040479063;
assign addr[42390]= 2015345591;
assign addr[42391]= 1987655498;
assign addr[42392]= 1957443913;
assign addr[42393]= 1924749160;
assign addr[42394]= 1889612716;
assign addr[42395]= 1852079154;
assign addr[42396]= 1812196087;
assign addr[42397]= 1770014111;
assign addr[42398]= 1725586737;
assign addr[42399]= 1678970324;
assign addr[42400]= 1630224009;
assign addr[42401]= 1579409630;
assign addr[42402]= 1526591649;
assign addr[42403]= 1471837070;
assign addr[42404]= 1415215352;
assign addr[42405]= 1356798326;
assign addr[42406]= 1296660098;
assign addr[42407]= 1234876957;
assign addr[42408]= 1171527280;
assign addr[42409]= 1106691431;
assign addr[42410]= 1040451659;
assign addr[42411]= 972891995;
assign addr[42412]= 904098143;
assign addr[42413]= 834157373;
assign addr[42414]= 763158411;
assign addr[42415]= 691191324;
assign addr[42416]= 618347408;
assign addr[42417]= 544719071;
assign addr[42418]= 470399716;
assign addr[42419]= 395483624;
assign addr[42420]= 320065829;
assign addr[42421]= 244242007;
assign addr[42422]= 168108346;
assign addr[42423]= 91761426;
assign addr[42424]= 15298099;
assign addr[42425]= -61184634;
assign addr[42426]= -137589750;
assign addr[42427]= -213820322;
assign addr[42428]= -289779648;
assign addr[42429]= -365371365;
assign addr[42430]= -440499581;
assign addr[42431]= -515068990;
assign addr[42432]= -588984994;
assign addr[42433]= -662153826;
assign addr[42434]= -734482665;
assign addr[42435]= -805879757;
assign addr[42436]= -876254528;
assign addr[42437]= -945517704;
assign addr[42438]= -1013581418;
assign addr[42439]= -1080359326;
assign addr[42440]= -1145766716;
assign addr[42441]= -1209720613;
assign addr[42442]= -1272139887;
assign addr[42443]= -1332945355;
assign addr[42444]= -1392059879;
assign addr[42445]= -1449408469;
assign addr[42446]= -1504918373;
assign addr[42447]= -1558519173;
assign addr[42448]= -1610142873;
assign addr[42449]= -1659723983;
assign addr[42450]= -1707199606;
assign addr[42451]= -1752509516;
assign addr[42452]= -1795596234;
assign addr[42453]= -1836405100;
assign addr[42454]= -1874884346;
assign addr[42455]= -1910985158;
assign addr[42456]= -1944661739;
assign addr[42457]= -1975871368;
assign addr[42458]= -2004574453;
assign addr[42459]= -2030734582;
assign addr[42460]= -2054318569;
assign addr[42461]= -2075296495;
assign addr[42462]= -2093641749;
assign addr[42463]= -2109331059;
assign addr[42464]= -2122344521;
assign addr[42465]= -2132665626;
assign addr[42466]= -2140281282;
assign addr[42467]= -2145181827;
assign addr[42468]= -2147361045;
assign addr[42469]= -2146816171;
assign addr[42470]= -2143547897;
assign addr[42471]= -2137560369;
assign addr[42472]= -2128861181;
assign addr[42473]= -2117461370;
assign addr[42474]= -2103375398;
assign addr[42475]= -2086621133;
assign addr[42476]= -2067219829;
assign addr[42477]= -2045196100;
assign addr[42478]= -2020577882;
assign addr[42479]= -1993396407;
assign addr[42480]= -1963686155;
assign addr[42481]= -1931484818;
assign addr[42482]= -1896833245;
assign addr[42483]= -1859775393;
assign addr[42484]= -1820358275;
assign addr[42485]= -1778631892;
assign addr[42486]= -1734649179;
assign addr[42487]= -1688465931;
assign addr[42488]= -1640140734;
assign addr[42489]= -1589734894;
assign addr[42490]= -1537312353;
assign addr[42491]= -1482939614;
assign addr[42492]= -1426685652;
assign addr[42493]= -1368621831;
assign addr[42494]= -1308821808;
assign addr[42495]= -1247361445;
assign addr[42496]= -1184318708;
assign addr[42497]= -1119773573;
assign addr[42498]= -1053807919;
assign addr[42499]= -986505429;
assign addr[42500]= -917951481;
assign addr[42501]= -848233042;
assign addr[42502]= -777438554;
assign addr[42503]= -705657826;
assign addr[42504]= -632981917;
assign addr[42505]= -559503022;
assign addr[42506]= -485314355;
assign addr[42507]= -410510029;
assign addr[42508]= -335184940;
assign addr[42509]= -259434643;
assign addr[42510]= -183355234;
assign addr[42511]= -107043224;
assign addr[42512]= -30595422;
assign addr[42513]= 45891193;
assign addr[42514]= 122319591;
assign addr[42515]= 198592817;
assign addr[42516]= 274614114;
assign addr[42517]= 350287041;
assign addr[42518]= 425515602;
assign addr[42519]= 500204365;
assign addr[42520]= 574258580;
assign addr[42521]= 647584304;
assign addr[42522]= 720088517;
assign addr[42523]= 791679244;
assign addr[42524]= 862265664;
assign addr[42525]= 931758235;
assign addr[42526]= 1000068799;
assign addr[42527]= 1067110699;
assign addr[42528]= 1132798888;
assign addr[42529]= 1197050035;
assign addr[42530]= 1259782632;
assign addr[42531]= 1320917099;
assign addr[42532]= 1380375881;
assign addr[42533]= 1438083551;
assign addr[42534]= 1493966902;
assign addr[42535]= 1547955041;
assign addr[42536]= 1599979481;
assign addr[42537]= 1649974225;
assign addr[42538]= 1697875851;
assign addr[42539]= 1743623590;
assign addr[42540]= 1787159411;
assign addr[42541]= 1828428082;
assign addr[42542]= 1867377253;
assign addr[42543]= 1903957513;
assign addr[42544]= 1938122457;
assign addr[42545]= 1969828744;
assign addr[42546]= 1999036154;
assign addr[42547]= 2025707632;
assign addr[42548]= 2049809346;
assign addr[42549]= 2071310720;
assign addr[42550]= 2090184478;
assign addr[42551]= 2106406677;
assign addr[42552]= 2119956737;
assign addr[42553]= 2130817471;
assign addr[42554]= 2138975100;
assign addr[42555]= 2144419275;
assign addr[42556]= 2147143090;
assign addr[42557]= 2147143090;
assign addr[42558]= 2144419275;
assign addr[42559]= 2138975100;
assign addr[42560]= 2130817471;
assign addr[42561]= 2119956737;
assign addr[42562]= 2106406677;
assign addr[42563]= 2090184478;
assign addr[42564]= 2071310720;
assign addr[42565]= 2049809346;
assign addr[42566]= 2025707632;
assign addr[42567]= 1999036154;
assign addr[42568]= 1969828744;
assign addr[42569]= 1938122457;
assign addr[42570]= 1903957513;
assign addr[42571]= 1867377253;
assign addr[42572]= 1828428082;
assign addr[42573]= 1787159411;
assign addr[42574]= 1743623590;
assign addr[42575]= 1697875851;
assign addr[42576]= 1649974225;
assign addr[42577]= 1599979481;
assign addr[42578]= 1547955041;
assign addr[42579]= 1493966902;
assign addr[42580]= 1438083551;
assign addr[42581]= 1380375881;
assign addr[42582]= 1320917099;
assign addr[42583]= 1259782632;
assign addr[42584]= 1197050035;
assign addr[42585]= 1132798888;
assign addr[42586]= 1067110699;
assign addr[42587]= 1000068799;
assign addr[42588]= 931758235;
assign addr[42589]= 862265664;
assign addr[42590]= 791679244;
assign addr[42591]= 720088517;
assign addr[42592]= 647584304;
assign addr[42593]= 574258580;
assign addr[42594]= 500204365;
assign addr[42595]= 425515602;
assign addr[42596]= 350287041;
assign addr[42597]= 274614114;
assign addr[42598]= 198592817;
assign addr[42599]= 122319591;
assign addr[42600]= 45891193;
assign addr[42601]= -30595422;
assign addr[42602]= -107043224;
assign addr[42603]= -183355234;
assign addr[42604]= -259434643;
assign addr[42605]= -335184940;
assign addr[42606]= -410510029;
assign addr[42607]= -485314355;
assign addr[42608]= -559503022;
assign addr[42609]= -632981917;
assign addr[42610]= -705657826;
assign addr[42611]= -777438554;
assign addr[42612]= -848233042;
assign addr[42613]= -917951481;
assign addr[42614]= -986505429;
assign addr[42615]= -1053807919;
assign addr[42616]= -1119773573;
assign addr[42617]= -1184318708;
assign addr[42618]= -1247361445;
assign addr[42619]= -1308821808;
assign addr[42620]= -1368621831;
assign addr[42621]= -1426685652;
assign addr[42622]= -1482939614;
assign addr[42623]= -1537312353;
assign addr[42624]= -1589734894;
assign addr[42625]= -1640140734;
assign addr[42626]= -1688465931;
assign addr[42627]= -1734649179;
assign addr[42628]= -1778631892;
assign addr[42629]= -1820358275;
assign addr[42630]= -1859775393;
assign addr[42631]= -1896833245;
assign addr[42632]= -1931484818;
assign addr[42633]= -1963686155;
assign addr[42634]= -1993396407;
assign addr[42635]= -2020577882;
assign addr[42636]= -2045196100;
assign addr[42637]= -2067219829;
assign addr[42638]= -2086621133;
assign addr[42639]= -2103375398;
assign addr[42640]= -2117461370;
assign addr[42641]= -2128861181;
assign addr[42642]= -2137560369;
assign addr[42643]= -2143547897;
assign addr[42644]= -2146816171;
assign addr[42645]= -2147361045;
assign addr[42646]= -2145181827;
assign addr[42647]= -2140281282;
assign addr[42648]= -2132665626;
assign addr[42649]= -2122344521;
assign addr[42650]= -2109331059;
assign addr[42651]= -2093641749;
assign addr[42652]= -2075296495;
assign addr[42653]= -2054318569;
assign addr[42654]= -2030734582;
assign addr[42655]= -2004574453;
assign addr[42656]= -1975871368;
assign addr[42657]= -1944661739;
assign addr[42658]= -1910985158;
assign addr[42659]= -1874884346;
assign addr[42660]= -1836405100;
assign addr[42661]= -1795596234;
assign addr[42662]= -1752509516;
assign addr[42663]= -1707199606;
assign addr[42664]= -1659723983;
assign addr[42665]= -1610142873;
assign addr[42666]= -1558519173;
assign addr[42667]= -1504918373;
assign addr[42668]= -1449408469;
assign addr[42669]= -1392059879;
assign addr[42670]= -1332945355;
assign addr[42671]= -1272139887;
assign addr[42672]= -1209720613;
assign addr[42673]= -1145766716;
assign addr[42674]= -1080359326;
assign addr[42675]= -1013581418;
assign addr[42676]= -945517704;
assign addr[42677]= -876254528;
assign addr[42678]= -805879757;
assign addr[42679]= -734482665;
assign addr[42680]= -662153826;
assign addr[42681]= -588984994;
assign addr[42682]= -515068990;
assign addr[42683]= -440499581;
assign addr[42684]= -365371365;
assign addr[42685]= -289779648;
assign addr[42686]= -213820322;
assign addr[42687]= -137589750;
assign addr[42688]= -61184634;
assign addr[42689]= 15298099;
assign addr[42690]= 91761426;
assign addr[42691]= 168108346;
assign addr[42692]= 244242007;
assign addr[42693]= 320065829;
assign addr[42694]= 395483624;
assign addr[42695]= 470399716;
assign addr[42696]= 544719071;
assign addr[42697]= 618347408;
assign addr[42698]= 691191324;
assign addr[42699]= 763158411;
assign addr[42700]= 834157373;
assign addr[42701]= 904098143;
assign addr[42702]= 972891995;
assign addr[42703]= 1040451659;
assign addr[42704]= 1106691431;
assign addr[42705]= 1171527280;
assign addr[42706]= 1234876957;
assign addr[42707]= 1296660098;
assign addr[42708]= 1356798326;
assign addr[42709]= 1415215352;
assign addr[42710]= 1471837070;
assign addr[42711]= 1526591649;
assign addr[42712]= 1579409630;
assign addr[42713]= 1630224009;
assign addr[42714]= 1678970324;
assign addr[42715]= 1725586737;
assign addr[42716]= 1770014111;
assign addr[42717]= 1812196087;
assign addr[42718]= 1852079154;
assign addr[42719]= 1889612716;
assign addr[42720]= 1924749160;
assign addr[42721]= 1957443913;
assign addr[42722]= 1987655498;
assign addr[42723]= 2015345591;
assign addr[42724]= 2040479063;
assign addr[42725]= 2063024031;
assign addr[42726]= 2082951896;
assign addr[42727]= 2100237377;
assign addr[42728]= 2114858546;
assign addr[42729]= 2126796855;
assign addr[42730]= 2136037160;
assign addr[42731]= 2142567738;
assign addr[42732]= 2146380306;
assign addr[42733]= 2147470025;
assign addr[42734]= 2145835515;
assign addr[42735]= 2141478848;
assign addr[42736]= 2134405552;
assign addr[42737]= 2124624598;
assign addr[42738]= 2112148396;
assign addr[42739]= 2096992772;
assign addr[42740]= 2079176953;
assign addr[42741]= 2058723538;
assign addr[42742]= 2035658475;
assign addr[42743]= 2010011024;
assign addr[42744]= 1981813720;
assign addr[42745]= 1951102334;
assign addr[42746]= 1917915825;
assign addr[42747]= 1882296293;
assign addr[42748]= 1844288924;
assign addr[42749]= 1803941934;
assign addr[42750]= 1761306505;
assign addr[42751]= 1716436725;
assign addr[42752]= 1669389513;
assign addr[42753]= 1620224553;
assign addr[42754]= 1569004214;
assign addr[42755]= 1515793473;
assign addr[42756]= 1460659832;
assign addr[42757]= 1403673233;
assign addr[42758]= 1344905966;
assign addr[42759]= 1284432584;
assign addr[42760]= 1222329801;
assign addr[42761]= 1158676398;
assign addr[42762]= 1093553126;
assign addr[42763]= 1027042599;
assign addr[42764]= 959229189;
assign addr[42765]= 890198924;
assign addr[42766]= 820039373;
assign addr[42767]= 748839539;
assign addr[42768]= 676689746;
assign addr[42769]= 603681519;
assign addr[42770]= 529907477;
assign addr[42771]= 455461206;
assign addr[42772]= 380437148;
assign addr[42773]= 304930476;
assign addr[42774]= 229036977;
assign addr[42775]= 152852926;
assign addr[42776]= 76474970;
assign addr[42777]= 0;
assign addr[42778]= -76474970;
assign addr[42779]= -152852926;
assign addr[42780]= -229036977;
assign addr[42781]= -304930476;
assign addr[42782]= -380437148;
assign addr[42783]= -455461206;
assign addr[42784]= -529907477;
assign addr[42785]= -603681519;
assign addr[42786]= -676689746;
assign addr[42787]= -748839539;
assign addr[42788]= -820039373;
assign addr[42789]= -890198924;
assign addr[42790]= -959229189;
assign addr[42791]= -1027042599;
assign addr[42792]= -1093553126;
assign addr[42793]= -1158676398;
assign addr[42794]= -1222329801;
assign addr[42795]= -1284432584;
assign addr[42796]= -1344905966;
assign addr[42797]= -1403673233;
assign addr[42798]= -1460659832;
assign addr[42799]= -1515793473;
assign addr[42800]= -1569004214;
assign addr[42801]= -1620224553;
assign addr[42802]= -1669389513;
assign addr[42803]= -1716436725;
assign addr[42804]= -1761306505;
assign addr[42805]= -1803941934;
assign addr[42806]= -1844288924;
assign addr[42807]= -1882296293;
assign addr[42808]= -1917915825;
assign addr[42809]= -1951102334;
assign addr[42810]= -1981813720;
assign addr[42811]= -2010011024;
assign addr[42812]= -2035658475;
assign addr[42813]= -2058723538;
assign addr[42814]= -2079176953;
assign addr[42815]= -2096992772;
assign addr[42816]= -2112148396;
assign addr[42817]= -2124624598;
assign addr[42818]= -2134405552;
assign addr[42819]= -2141478848;
assign addr[42820]= -2145835515;
assign addr[42821]= -2147470025;
assign addr[42822]= -2146380306;
assign addr[42823]= -2142567738;
assign addr[42824]= -2136037160;
assign addr[42825]= -2126796855;
assign addr[42826]= -2114858546;
assign addr[42827]= -2100237377;
assign addr[42828]= -2082951896;
assign addr[42829]= -2063024031;
assign addr[42830]= -2040479063;
assign addr[42831]= -2015345591;
assign addr[42832]= -1987655498;
assign addr[42833]= -1957443913;
assign addr[42834]= -1924749160;
assign addr[42835]= -1889612716;
assign addr[42836]= -1852079154;
assign addr[42837]= -1812196087;
assign addr[42838]= -1770014111;
assign addr[42839]= -1725586737;
assign addr[42840]= -1678970324;
assign addr[42841]= -1630224009;
assign addr[42842]= -1579409630;
assign addr[42843]= -1526591649;
assign addr[42844]= -1471837070;
assign addr[42845]= -1415215352;
assign addr[42846]= -1356798326;
assign addr[42847]= -1296660098;
assign addr[42848]= -1234876957;
assign addr[42849]= -1171527280;
assign addr[42850]= -1106691431;
assign addr[42851]= -1040451659;
assign addr[42852]= -972891995;
assign addr[42853]= -904098143;
assign addr[42854]= -834157373;
assign addr[42855]= -763158411;
assign addr[42856]= -691191324;
assign addr[42857]= -618347408;
assign addr[42858]= -544719071;
assign addr[42859]= -470399716;
assign addr[42860]= -395483624;
assign addr[42861]= -320065829;
assign addr[42862]= -244242007;
assign addr[42863]= -168108346;
assign addr[42864]= -91761426;
assign addr[42865]= -15298099;
assign addr[42866]= 61184634;
assign addr[42867]= 137589750;
assign addr[42868]= 213820322;
assign addr[42869]= 289779648;
assign addr[42870]= 365371365;
assign addr[42871]= 440499581;
assign addr[42872]= 515068990;
assign addr[42873]= 588984994;
assign addr[42874]= 662153826;
assign addr[42875]= 734482665;
assign addr[42876]= 805879757;
assign addr[42877]= 876254528;
assign addr[42878]= 945517704;
assign addr[42879]= 1013581418;
assign addr[42880]= 1080359326;
assign addr[42881]= 1145766716;
assign addr[42882]= 1209720613;
assign addr[42883]= 1272139887;
assign addr[42884]= 1332945355;
assign addr[42885]= 1392059879;
assign addr[42886]= 1449408469;
assign addr[42887]= 1504918373;
assign addr[42888]= 1558519173;
assign addr[42889]= 1610142873;
assign addr[42890]= 1659723983;
assign addr[42891]= 1707199606;
assign addr[42892]= 1752509516;
assign addr[42893]= 1795596234;
assign addr[42894]= 1836405100;
assign addr[42895]= 1874884346;
assign addr[42896]= 1910985158;
assign addr[42897]= 1944661739;
assign addr[42898]= 1975871368;
assign addr[42899]= 2004574453;
assign addr[42900]= 2030734582;
assign addr[42901]= 2054318569;
assign addr[42902]= 2075296495;
assign addr[42903]= 2093641749;
assign addr[42904]= 2109331059;
assign addr[42905]= 2122344521;
assign addr[42906]= 2132665626;
assign addr[42907]= 2140281282;
assign addr[42908]= 2145181827;
assign addr[42909]= 2147361045;
assign addr[42910]= 2146816171;
assign addr[42911]= 2143547897;
assign addr[42912]= 2137560369;
assign addr[42913]= 2128861181;
assign addr[42914]= 2117461370;
assign addr[42915]= 2103375398;
assign addr[42916]= 2086621133;
assign addr[42917]= 2067219829;
assign addr[42918]= 2045196100;
assign addr[42919]= 2020577882;
assign addr[42920]= 1993396407;
assign addr[42921]= 1963686155;
assign addr[42922]= 1931484818;
assign addr[42923]= 1896833245;
assign addr[42924]= 1859775393;
assign addr[42925]= 1820358275;
assign addr[42926]= 1778631892;
assign addr[42927]= 1734649179;
assign addr[42928]= 1688465931;
assign addr[42929]= 1640140734;
assign addr[42930]= 1589734894;
assign addr[42931]= 1537312353;
assign addr[42932]= 1482939614;
assign addr[42933]= 1426685652;
assign addr[42934]= 1368621831;
assign addr[42935]= 1308821808;
assign addr[42936]= 1247361445;
assign addr[42937]= 1184318708;
assign addr[42938]= 1119773573;
assign addr[42939]= 1053807919;
assign addr[42940]= 986505429;
assign addr[42941]= 917951481;
assign addr[42942]= 848233042;
assign addr[42943]= 777438554;
assign addr[42944]= 705657826;
assign addr[42945]= 632981917;
assign addr[42946]= 559503022;
assign addr[42947]= 485314355;
assign addr[42948]= 410510029;
assign addr[42949]= 335184940;
assign addr[42950]= 259434643;
assign addr[42951]= 183355234;
assign addr[42952]= 107043224;
assign addr[42953]= 30595422;
assign addr[42954]= -45891193;
assign addr[42955]= -122319591;
assign addr[42956]= -198592817;
assign addr[42957]= -274614114;
assign addr[42958]= -350287041;
assign addr[42959]= -425515602;
assign addr[42960]= -500204365;
assign addr[42961]= -574258580;
assign addr[42962]= -647584304;
assign addr[42963]= -720088517;
assign addr[42964]= -791679244;
assign addr[42965]= -862265664;
assign addr[42966]= -931758235;
assign addr[42967]= -1000068799;
assign addr[42968]= -1067110699;
assign addr[42969]= -1132798888;
assign addr[42970]= -1197050035;
assign addr[42971]= -1259782632;
assign addr[42972]= -1320917099;
assign addr[42973]= -1380375881;
assign addr[42974]= -1438083551;
assign addr[42975]= -1493966902;
assign addr[42976]= -1547955041;
assign addr[42977]= -1599979481;
assign addr[42978]= -1649974225;
assign addr[42979]= -1697875851;
assign addr[42980]= -1743623590;
assign addr[42981]= -1787159411;
assign addr[42982]= -1828428082;
assign addr[42983]= -1867377253;
assign addr[42984]= -1903957513;
assign addr[42985]= -1938122457;
assign addr[42986]= -1969828744;
assign addr[42987]= -1999036154;
assign addr[42988]= -2025707632;
assign addr[42989]= -2049809346;
assign addr[42990]= -2071310720;
assign addr[42991]= -2090184478;
assign addr[42992]= -2106406677;
assign addr[42993]= -2119956737;
assign addr[42994]= -2130817471;
assign addr[42995]= -2138975100;
assign addr[42996]= -2144419275;
assign addr[42997]= -2147143090;
assign addr[42998]= -2147143090;
assign addr[42999]= -2144419275;
assign addr[43000]= -2138975100;
assign addr[43001]= -2130817471;
assign addr[43002]= -2119956737;
assign addr[43003]= -2106406677;
assign addr[43004]= -2090184478;
assign addr[43005]= -2071310720;
assign addr[43006]= -2049809346;
assign addr[43007]= -2025707632;
assign addr[43008]= -1999036154;
assign addr[43009]= -1969828744;
assign addr[43010]= -1938122457;
assign addr[43011]= -1903957513;
assign addr[43012]= -1867377253;
assign addr[43013]= -1828428082;
assign addr[43014]= -1787159411;
assign addr[43015]= -1743623590;
assign addr[43016]= -1697875851;
assign addr[43017]= -1649974225;
assign addr[43018]= -1599979481;
assign addr[43019]= -1547955041;
assign addr[43020]= -1493966902;
assign addr[43021]= -1438083551;
assign addr[43022]= -1380375881;
assign addr[43023]= -1320917099;
assign addr[43024]= -1259782632;
assign addr[43025]= -1197050035;
assign addr[43026]= -1132798888;
assign addr[43027]= -1067110699;
assign addr[43028]= -1000068799;
assign addr[43029]= -931758235;
assign addr[43030]= -862265664;
assign addr[43031]= -791679244;
assign addr[43032]= -720088517;
assign addr[43033]= -647584304;
assign addr[43034]= -574258580;
assign addr[43035]= -500204365;
assign addr[43036]= -425515602;
assign addr[43037]= -350287041;
assign addr[43038]= -274614114;
assign addr[43039]= -198592817;
assign addr[43040]= -122319591;
assign addr[43041]= -45891193;
assign addr[43042]= 30595422;
assign addr[43043]= 107043224;
assign addr[43044]= 183355234;
assign addr[43045]= 259434643;
assign addr[43046]= 335184940;
assign addr[43047]= 410510029;
assign addr[43048]= 485314355;
assign addr[43049]= 559503022;
assign addr[43050]= 632981917;
assign addr[43051]= 705657826;
assign addr[43052]= 777438554;
assign addr[43053]= 848233042;
assign addr[43054]= 917951481;
assign addr[43055]= 986505429;
assign addr[43056]= 1053807919;
assign addr[43057]= 1119773573;
assign addr[43058]= 1184318708;
assign addr[43059]= 1247361445;
assign addr[43060]= 1308821808;
assign addr[43061]= 1368621831;
assign addr[43062]= 1426685652;
assign addr[43063]= 1482939614;
assign addr[43064]= 1537312353;
assign addr[43065]= 1589734894;
assign addr[43066]= 1640140734;
assign addr[43067]= 1688465931;
assign addr[43068]= 1734649179;
assign addr[43069]= 1778631892;
assign addr[43070]= 1820358275;
assign addr[43071]= 1859775393;
assign addr[43072]= 1896833245;
assign addr[43073]= 1931484818;
assign addr[43074]= 1963686155;
assign addr[43075]= 1993396407;
assign addr[43076]= 2020577882;
assign addr[43077]= 2045196100;
assign addr[43078]= 2067219829;
assign addr[43079]= 2086621133;
assign addr[43080]= 2103375398;
assign addr[43081]= 2117461370;
assign addr[43082]= 2128861181;
assign addr[43083]= 2137560369;
assign addr[43084]= 2143547897;
assign addr[43085]= 2146816171;
assign addr[43086]= 2147361045;
assign addr[43087]= 2145181827;
assign addr[43088]= 2140281282;
assign addr[43089]= 2132665626;
assign addr[43090]= 2122344521;
assign addr[43091]= 2109331059;
assign addr[43092]= 2093641749;
assign addr[43093]= 2075296495;
assign addr[43094]= 2054318569;
assign addr[43095]= 2030734582;
assign addr[43096]= 2004574453;
assign addr[43097]= 1975871368;
assign addr[43098]= 1944661739;
assign addr[43099]= 1910985158;
assign addr[43100]= 1874884346;
assign addr[43101]= 1836405100;
assign addr[43102]= 1795596234;
assign addr[43103]= 1752509516;
assign addr[43104]= 1707199606;
assign addr[43105]= 1659723983;
assign addr[43106]= 1610142873;
assign addr[43107]= 1558519173;
assign addr[43108]= 1504918373;
assign addr[43109]= 1449408469;
assign addr[43110]= 1392059879;
assign addr[43111]= 1332945355;
assign addr[43112]= 1272139887;
assign addr[43113]= 1209720613;
assign addr[43114]= 1145766716;
assign addr[43115]= 1080359326;
assign addr[43116]= 1013581418;
assign addr[43117]= 945517704;
assign addr[43118]= 876254528;
assign addr[43119]= 805879757;
assign addr[43120]= 734482665;
assign addr[43121]= 662153826;
assign addr[43122]= 588984994;
assign addr[43123]= 515068990;
assign addr[43124]= 440499581;
assign addr[43125]= 365371365;
assign addr[43126]= 289779648;
assign addr[43127]= 213820322;
assign addr[43128]= 137589750;
assign addr[43129]= 61184634;
assign addr[43130]= -15298099;
assign addr[43131]= -91761426;
assign addr[43132]= -168108346;
assign addr[43133]= -244242007;
assign addr[43134]= -320065829;
assign addr[43135]= -395483624;
assign addr[43136]= -470399716;
assign addr[43137]= -544719071;
assign addr[43138]= -618347408;
assign addr[43139]= -691191324;
assign addr[43140]= -763158411;
assign addr[43141]= -834157373;
assign addr[43142]= -904098143;
assign addr[43143]= -972891995;
assign addr[43144]= -1040451659;
assign addr[43145]= -1106691431;
assign addr[43146]= -1171527280;
assign addr[43147]= -1234876957;
assign addr[43148]= -1296660098;
assign addr[43149]= -1356798326;
assign addr[43150]= -1415215352;
assign addr[43151]= -1471837070;
assign addr[43152]= -1526591649;
assign addr[43153]= -1579409630;
assign addr[43154]= -1630224009;
assign addr[43155]= -1678970324;
assign addr[43156]= -1725586737;
assign addr[43157]= -1770014111;
assign addr[43158]= -1812196087;
assign addr[43159]= -1852079154;
assign addr[43160]= -1889612716;
assign addr[43161]= -1924749160;
assign addr[43162]= -1957443913;
assign addr[43163]= -1987655498;
assign addr[43164]= -2015345591;
assign addr[43165]= -2040479063;
assign addr[43166]= -2063024031;
assign addr[43167]= -2082951896;
assign addr[43168]= -2100237377;
assign addr[43169]= -2114858546;
assign addr[43170]= -2126796855;
assign addr[43171]= -2136037160;
assign addr[43172]= -2142567738;
assign addr[43173]= -2146380306;
assign addr[43174]= -2147470025;
assign addr[43175]= -2145835515;
assign addr[43176]= -2141478848;
assign addr[43177]= -2134405552;
assign addr[43178]= -2124624598;
assign addr[43179]= -2112148396;
assign addr[43180]= -2096992772;
assign addr[43181]= -2079176953;
assign addr[43182]= -2058723538;
assign addr[43183]= -2035658475;
assign addr[43184]= -2010011024;
assign addr[43185]= -1981813720;
assign addr[43186]= -1951102334;
assign addr[43187]= -1917915825;
assign addr[43188]= -1882296293;
assign addr[43189]= -1844288924;
assign addr[43190]= -1803941934;
assign addr[43191]= -1761306505;
assign addr[43192]= -1716436725;
assign addr[43193]= -1669389513;
assign addr[43194]= -1620224553;
assign addr[43195]= -1569004214;
assign addr[43196]= -1515793473;
assign addr[43197]= -1460659832;
assign addr[43198]= -1403673233;
assign addr[43199]= -1344905966;
assign addr[43200]= -1284432584;
assign addr[43201]= -1222329801;
assign addr[43202]= -1158676398;
assign addr[43203]= -1093553126;
assign addr[43204]= -1027042599;
assign addr[43205]= -959229189;
assign addr[43206]= -890198924;
assign addr[43207]= -820039373;
assign addr[43208]= -748839539;
assign addr[43209]= -676689746;
assign addr[43210]= -603681519;
assign addr[43211]= -529907477;
assign addr[43212]= -455461206;
assign addr[43213]= -380437148;
assign addr[43214]= -304930476;
assign addr[43215]= -229036977;
assign addr[43216]= -152852926;
assign addr[43217]= -76474970;
assign addr[43218]= 0;
assign addr[43219]= 76474970;
assign addr[43220]= 152852926;
assign addr[43221]= 229036977;
assign addr[43222]= 304930476;
assign addr[43223]= 380437148;
assign addr[43224]= 455461206;
assign addr[43225]= 529907477;
assign addr[43226]= 603681519;
assign addr[43227]= 676689746;
assign addr[43228]= 748839539;
assign addr[43229]= 820039373;
assign addr[43230]= 890198924;
assign addr[43231]= 959229189;
assign addr[43232]= 1027042599;
assign addr[43233]= 1093553126;
assign addr[43234]= 1158676398;
assign addr[43235]= 1222329801;
assign addr[43236]= 1284432584;
assign addr[43237]= 1344905966;
assign addr[43238]= 1403673233;
assign addr[43239]= 1460659832;
assign addr[43240]= 1515793473;
assign addr[43241]= 1569004214;
assign addr[43242]= 1620224553;
assign addr[43243]= 1669389513;
assign addr[43244]= 1716436725;
assign addr[43245]= 1761306505;
assign addr[43246]= 1803941934;
assign addr[43247]= 1844288924;
assign addr[43248]= 1882296293;
assign addr[43249]= 1917915825;
assign addr[43250]= 1951102334;
assign addr[43251]= 1981813720;
assign addr[43252]= 2010011024;
assign addr[43253]= 2035658475;
assign addr[43254]= 2058723538;
assign addr[43255]= 2079176953;
assign addr[43256]= 2096992772;
assign addr[43257]= 2112148396;
assign addr[43258]= 2124624598;
assign addr[43259]= 2134405552;
assign addr[43260]= 2141478848;
assign addr[43261]= 2145835515;
assign addr[43262]= 2147470025;
assign addr[43263]= 2146380306;
assign addr[43264]= 2142567738;
assign addr[43265]= 2136037160;
assign addr[43266]= 2126796855;
assign addr[43267]= 2114858546;
assign addr[43268]= 2100237377;
assign addr[43269]= 2082951896;
assign addr[43270]= 2063024031;
assign addr[43271]= 2040479063;
assign addr[43272]= 2015345591;
assign addr[43273]= 1987655498;
assign addr[43274]= 1957443913;
assign addr[43275]= 1924749160;
assign addr[43276]= 1889612716;
assign addr[43277]= 1852079154;
assign addr[43278]= 1812196087;
assign addr[43279]= 1770014111;
assign addr[43280]= 1725586737;
assign addr[43281]= 1678970324;
assign addr[43282]= 1630224009;
assign addr[43283]= 1579409630;
assign addr[43284]= 1526591649;
assign addr[43285]= 1471837070;
assign addr[43286]= 1415215352;
assign addr[43287]= 1356798326;
assign addr[43288]= 1296660098;
assign addr[43289]= 1234876957;
assign addr[43290]= 1171527280;
assign addr[43291]= 1106691431;
assign addr[43292]= 1040451659;
assign addr[43293]= 972891995;
assign addr[43294]= 904098143;
assign addr[43295]= 834157373;
assign addr[43296]= 763158411;
assign addr[43297]= 691191324;
assign addr[43298]= 618347408;
assign addr[43299]= 544719071;
assign addr[43300]= 470399716;
assign addr[43301]= 395483624;
assign addr[43302]= 320065829;
assign addr[43303]= 244242007;
assign addr[43304]= 168108346;
assign addr[43305]= 91761426;
assign addr[43306]= 15298099;
assign addr[43307]= -61184634;
assign addr[43308]= -137589750;
assign addr[43309]= -213820322;
assign addr[43310]= -289779648;
assign addr[43311]= -365371365;
assign addr[43312]= -440499581;
assign addr[43313]= -515068990;
assign addr[43314]= -588984994;
assign addr[43315]= -662153826;
assign addr[43316]= -734482665;
assign addr[43317]= -805879757;
assign addr[43318]= -876254528;
assign addr[43319]= -945517704;
assign addr[43320]= -1013581418;
assign addr[43321]= -1080359326;
assign addr[43322]= -1145766716;
assign addr[43323]= -1209720613;
assign addr[43324]= -1272139887;
assign addr[43325]= -1332945355;
assign addr[43326]= -1392059879;
assign addr[43327]= -1449408469;
assign addr[43328]= -1504918373;
assign addr[43329]= -1558519173;
assign addr[43330]= -1610142873;
assign addr[43331]= -1659723983;
assign addr[43332]= -1707199606;
assign addr[43333]= -1752509516;
assign addr[43334]= -1795596234;
assign addr[43335]= -1836405100;
assign addr[43336]= -1874884346;
assign addr[43337]= -1910985158;
assign addr[43338]= -1944661739;
assign addr[43339]= -1975871368;
assign addr[43340]= -2004574453;
assign addr[43341]= -2030734582;
assign addr[43342]= -2054318569;
assign addr[43343]= -2075296495;
assign addr[43344]= -2093641749;
assign addr[43345]= -2109331059;
assign addr[43346]= -2122344521;
assign addr[43347]= -2132665626;
assign addr[43348]= -2140281282;
assign addr[43349]= -2145181827;
assign addr[43350]= -2147361045;
assign addr[43351]= -2146816171;
assign addr[43352]= -2143547897;
assign addr[43353]= -2137560369;
assign addr[43354]= -2128861181;
assign addr[43355]= -2117461370;
assign addr[43356]= -2103375398;
assign addr[43357]= -2086621133;
assign addr[43358]= -2067219829;
assign addr[43359]= -2045196100;
assign addr[43360]= -2020577882;
assign addr[43361]= -1993396407;
assign addr[43362]= -1963686155;
assign addr[43363]= -1931484818;
assign addr[43364]= -1896833245;
assign addr[43365]= -1859775393;
assign addr[43366]= -1820358275;
assign addr[43367]= -1778631892;
assign addr[43368]= -1734649179;
assign addr[43369]= -1688465931;
assign addr[43370]= -1640140734;
assign addr[43371]= -1589734894;
assign addr[43372]= -1537312353;
assign addr[43373]= -1482939614;
assign addr[43374]= -1426685652;
assign addr[43375]= -1368621831;
assign addr[43376]= -1308821808;
assign addr[43377]= -1247361445;
assign addr[43378]= -1184318708;
assign addr[43379]= -1119773573;
assign addr[43380]= -1053807919;
assign addr[43381]= -986505429;
assign addr[43382]= -917951481;
assign addr[43383]= -848233042;
assign addr[43384]= -777438554;
assign addr[43385]= -705657826;
assign addr[43386]= -632981917;
assign addr[43387]= -559503022;
assign addr[43388]= -485314355;
assign addr[43389]= -410510029;
assign addr[43390]= -335184940;
assign addr[43391]= -259434643;
assign addr[43392]= -183355234;
assign addr[43393]= -107043224;
assign addr[43394]= -30595422;
assign addr[43395]= 45891193;
assign addr[43396]= 122319591;
assign addr[43397]= 198592817;
assign addr[43398]= 274614114;
assign addr[43399]= 350287041;
assign addr[43400]= 425515602;
assign addr[43401]= 500204365;
assign addr[43402]= 574258580;
assign addr[43403]= 647584304;
assign addr[43404]= 720088517;
assign addr[43405]= 791679244;
assign addr[43406]= 862265664;
assign addr[43407]= 931758235;
assign addr[43408]= 1000068799;
assign addr[43409]= 1067110699;
assign addr[43410]= 1132798888;
assign addr[43411]= 1197050035;
assign addr[43412]= 1259782632;
assign addr[43413]= 1320917099;
assign addr[43414]= 1380375881;
assign addr[43415]= 1438083551;
assign addr[43416]= 1493966902;
assign addr[43417]= 1547955041;
assign addr[43418]= 1599979481;
assign addr[43419]= 1649974225;
assign addr[43420]= 1697875851;
assign addr[43421]= 1743623590;
assign addr[43422]= 1787159411;
assign addr[43423]= 1828428082;
assign addr[43424]= 1867377253;
assign addr[43425]= 1903957513;
assign addr[43426]= 1938122457;
assign addr[43427]= 1969828744;
assign addr[43428]= 1999036154;
assign addr[43429]= 2025707632;
assign addr[43430]= 2049809346;
assign addr[43431]= 2071310720;
assign addr[43432]= 2090184478;
assign addr[43433]= 2106406677;
assign addr[43434]= 2119956737;
assign addr[43435]= 2130817471;
assign addr[43436]= 2138975100;
assign addr[43437]= 2144419275;
assign addr[43438]= 2147143090;
assign addr[43439]= 2147143090;
assign addr[43440]= 2144419275;
assign addr[43441]= 2138975100;
assign addr[43442]= 2130817471;
assign addr[43443]= 2119956737;
assign addr[43444]= 2106406677;
assign addr[43445]= 2090184478;
assign addr[43446]= 2071310720;
assign addr[43447]= 2049809346;
assign addr[43448]= 2025707632;
assign addr[43449]= 1999036154;
assign addr[43450]= 1969828744;
assign addr[43451]= 1938122457;
assign addr[43452]= 1903957513;
assign addr[43453]= 1867377253;
assign addr[43454]= 1828428082;
assign addr[43455]= 1787159411;
assign addr[43456]= 1743623590;
assign addr[43457]= 1697875851;
assign addr[43458]= 1649974225;
assign addr[43459]= 1599979481;
assign addr[43460]= 1547955041;
assign addr[43461]= 1493966902;
assign addr[43462]= 1438083551;
assign addr[43463]= 1380375881;
assign addr[43464]= 1320917099;
assign addr[43465]= 1259782632;
assign addr[43466]= 1197050035;
assign addr[43467]= 1132798888;
assign addr[43468]= 1067110699;
assign addr[43469]= 1000068799;
assign addr[43470]= 931758235;
assign addr[43471]= 862265664;
assign addr[43472]= 791679244;
assign addr[43473]= 720088517;
assign addr[43474]= 647584304;
assign addr[43475]= 574258580;
assign addr[43476]= 500204365;
assign addr[43477]= 425515602;
assign addr[43478]= 350287041;
assign addr[43479]= 274614114;
assign addr[43480]= 198592817;
assign addr[43481]= 122319591;
assign addr[43482]= 45891193;
assign addr[43483]= -30595422;
assign addr[43484]= -107043224;
assign addr[43485]= -183355234;
assign addr[43486]= -259434643;
assign addr[43487]= -335184940;
assign addr[43488]= -410510029;
assign addr[43489]= -485314355;
assign addr[43490]= -559503022;
assign addr[43491]= -632981917;
assign addr[43492]= -705657826;
assign addr[43493]= -777438554;
assign addr[43494]= -848233042;
assign addr[43495]= -917951481;
assign addr[43496]= -986505429;
assign addr[43497]= -1053807919;
assign addr[43498]= -1119773573;
assign addr[43499]= -1184318708;
assign addr[43500]= -1247361445;
assign addr[43501]= -1308821808;
assign addr[43502]= -1368621831;
assign addr[43503]= -1426685652;
assign addr[43504]= -1482939614;
assign addr[43505]= -1537312353;
assign addr[43506]= -1589734894;
assign addr[43507]= -1640140734;
assign addr[43508]= -1688465931;
assign addr[43509]= -1734649179;
assign addr[43510]= -1778631892;
assign addr[43511]= -1820358275;
assign addr[43512]= -1859775393;
assign addr[43513]= -1896833245;
assign addr[43514]= -1931484818;
assign addr[43515]= -1963686155;
assign addr[43516]= -1993396407;
assign addr[43517]= -2020577882;
assign addr[43518]= -2045196100;
assign addr[43519]= -2067219829;
assign addr[43520]= -2086621133;
assign addr[43521]= -2103375398;
assign addr[43522]= -2117461370;
assign addr[43523]= -2128861181;
assign addr[43524]= -2137560369;
assign addr[43525]= -2143547897;
assign addr[43526]= -2146816171;
assign addr[43527]= -2147361045;
assign addr[43528]= -2145181827;
assign addr[43529]= -2140281282;
assign addr[43530]= -2132665626;
assign addr[43531]= -2122344521;
assign addr[43532]= -2109331059;
assign addr[43533]= -2093641749;
assign addr[43534]= -2075296495;
assign addr[43535]= -2054318569;
assign addr[43536]= -2030734582;
assign addr[43537]= -2004574453;
assign addr[43538]= -1975871368;
assign addr[43539]= -1944661739;
assign addr[43540]= -1910985158;
assign addr[43541]= -1874884346;
assign addr[43542]= -1836405100;
assign addr[43543]= -1795596234;
assign addr[43544]= -1752509516;
assign addr[43545]= -1707199606;
assign addr[43546]= -1659723983;
assign addr[43547]= -1610142873;
assign addr[43548]= -1558519173;
assign addr[43549]= -1504918373;
assign addr[43550]= -1449408469;
assign addr[43551]= -1392059879;
assign addr[43552]= -1332945355;
assign addr[43553]= -1272139887;
assign addr[43554]= -1209720613;
assign addr[43555]= -1145766716;
assign addr[43556]= -1080359326;
assign addr[43557]= -1013581418;
assign addr[43558]= -945517704;
assign addr[43559]= -876254528;
assign addr[43560]= -805879757;
assign addr[43561]= -734482665;
assign addr[43562]= -662153826;
assign addr[43563]= -588984994;
assign addr[43564]= -515068990;
assign addr[43565]= -440499581;
assign addr[43566]= -365371365;
assign addr[43567]= -289779648;
assign addr[43568]= -213820322;
assign addr[43569]= -137589750;
assign addr[43570]= -61184634;
assign addr[43571]= 15298099;
assign addr[43572]= 91761426;
assign addr[43573]= 168108346;
assign addr[43574]= 244242007;
assign addr[43575]= 320065829;
assign addr[43576]= 395483624;
assign addr[43577]= 470399716;
assign addr[43578]= 544719071;
assign addr[43579]= 618347408;
assign addr[43580]= 691191324;
assign addr[43581]= 763158411;
assign addr[43582]= 834157373;
assign addr[43583]= 904098143;
assign addr[43584]= 972891995;
assign addr[43585]= 1040451659;
assign addr[43586]= 1106691431;
assign addr[43587]= 1171527280;
assign addr[43588]= 1234876957;
assign addr[43589]= 1296660098;
assign addr[43590]= 1356798326;
assign addr[43591]= 1415215352;
assign addr[43592]= 1471837070;
assign addr[43593]= 1526591649;
assign addr[43594]= 1579409630;
assign addr[43595]= 1630224009;
assign addr[43596]= 1678970324;
assign addr[43597]= 1725586737;
assign addr[43598]= 1770014111;
assign addr[43599]= 1812196087;
assign addr[43600]= 1852079154;
assign addr[43601]= 1889612716;
assign addr[43602]= 1924749160;
assign addr[43603]= 1957443913;
assign addr[43604]= 1987655498;
assign addr[43605]= 2015345591;
assign addr[43606]= 2040479063;
assign addr[43607]= 2063024031;
assign addr[43608]= 2082951896;
assign addr[43609]= 2100237377;
assign addr[43610]= 2114858546;
assign addr[43611]= 2126796855;
assign addr[43612]= 2136037160;
assign addr[43613]= 2142567738;
assign addr[43614]= 2146380306;
assign addr[43615]= 2147470025;
assign addr[43616]= 2145835515;
assign addr[43617]= 2141478848;
assign addr[43618]= 2134405552;
assign addr[43619]= 2124624598;
assign addr[43620]= 2112148396;
assign addr[43621]= 2096992772;
assign addr[43622]= 2079176953;
assign addr[43623]= 2058723538;
assign addr[43624]= 2035658475;
assign addr[43625]= 2010011024;
assign addr[43626]= 1981813720;
assign addr[43627]= 1951102334;
assign addr[43628]= 1917915825;
assign addr[43629]= 1882296293;
assign addr[43630]= 1844288924;
assign addr[43631]= 1803941934;
assign addr[43632]= 1761306505;
assign addr[43633]= 1716436725;
assign addr[43634]= 1669389513;
assign addr[43635]= 1620224553;
assign addr[43636]= 1569004214;
assign addr[43637]= 1515793473;
assign addr[43638]= 1460659832;
assign addr[43639]= 1403673233;
assign addr[43640]= 1344905966;
assign addr[43641]= 1284432584;
assign addr[43642]= 1222329801;
assign addr[43643]= 1158676398;
assign addr[43644]= 1093553126;
assign addr[43645]= 1027042599;
assign addr[43646]= 959229189;
assign addr[43647]= 890198924;
assign addr[43648]= 820039373;
assign addr[43649]= 748839539;
assign addr[43650]= 676689746;
assign addr[43651]= 603681519;
assign addr[43652]= 529907477;
assign addr[43653]= 455461206;
assign addr[43654]= 380437148;
assign addr[43655]= 304930476;
assign addr[43656]= 229036977;
assign addr[43657]= 152852926;
assign addr[43658]= 76474970;
assign addr[43659]= 0;
assign addr[43660]= -76474970;
assign addr[43661]= -152852926;
assign addr[43662]= -229036977;
assign addr[43663]= -304930476;
assign addr[43664]= -380437148;
assign addr[43665]= -455461206;
assign addr[43666]= -529907477;
assign addr[43667]= -603681519;
assign addr[43668]= -676689746;
assign addr[43669]= -748839539;
assign addr[43670]= -820039373;
assign addr[43671]= -890198924;
assign addr[43672]= -959229189;
assign addr[43673]= -1027042599;
assign addr[43674]= -1093553126;
assign addr[43675]= -1158676398;
assign addr[43676]= -1222329801;
assign addr[43677]= -1284432584;
assign addr[43678]= -1344905966;
assign addr[43679]= -1403673233;
assign addr[43680]= -1460659832;
assign addr[43681]= -1515793473;
assign addr[43682]= -1569004214;
assign addr[43683]= -1620224553;
assign addr[43684]= -1669389513;
assign addr[43685]= -1716436725;
assign addr[43686]= -1761306505;
assign addr[43687]= -1803941934;
assign addr[43688]= -1844288924;
assign addr[43689]= -1882296293;
assign addr[43690]= -1917915825;
assign addr[43691]= -1951102334;
assign addr[43692]= -1981813720;
assign addr[43693]= -2010011024;
assign addr[43694]= -2035658475;
assign addr[43695]= -2058723538;
assign addr[43696]= -2079176953;
assign addr[43697]= -2096992772;
assign addr[43698]= -2112148396;
assign addr[43699]= -2124624598;
assign addr[43700]= -2134405552;
assign addr[43701]= -2141478848;
assign addr[43702]= -2145835515;
assign addr[43703]= -2147470025;
assign addr[43704]= -2146380306;
assign addr[43705]= -2142567738;
assign addr[43706]= -2136037160;
assign addr[43707]= -2126796855;
assign addr[43708]= -2114858546;
assign addr[43709]= -2100237377;
assign addr[43710]= -2082951896;
assign addr[43711]= -2063024031;
assign addr[43712]= -2040479063;
assign addr[43713]= -2015345591;
assign addr[43714]= -1987655498;
assign addr[43715]= -1957443913;
assign addr[43716]= -1924749160;
assign addr[43717]= -1889612716;
assign addr[43718]= -1852079154;
assign addr[43719]= -1812196087;
assign addr[43720]= -1770014111;
assign addr[43721]= -1725586737;
assign addr[43722]= -1678970324;
assign addr[43723]= -1630224009;
assign addr[43724]= -1579409630;
assign addr[43725]= -1526591649;
assign addr[43726]= -1471837070;
assign addr[43727]= -1415215352;
assign addr[43728]= -1356798326;
assign addr[43729]= -1296660098;
assign addr[43730]= -1234876957;
assign addr[43731]= -1171527280;
assign addr[43732]= -1106691431;
assign addr[43733]= -1040451659;
assign addr[43734]= -972891995;
assign addr[43735]= -904098143;
assign addr[43736]= -834157373;
assign addr[43737]= -763158411;
assign addr[43738]= -691191324;
assign addr[43739]= -618347408;
assign addr[43740]= -544719071;
assign addr[43741]= -470399716;
assign addr[43742]= -395483624;
assign addr[43743]= -320065829;
assign addr[43744]= -244242007;
assign addr[43745]= -168108346;
assign addr[43746]= -91761426;
assign addr[43747]= -15298099;
assign addr[43748]= 61184634;
assign addr[43749]= 137589750;
assign addr[43750]= 213820322;
assign addr[43751]= 289779648;
assign addr[43752]= 365371365;
assign addr[43753]= 440499581;
assign addr[43754]= 515068990;
assign addr[43755]= 588984994;
assign addr[43756]= 662153826;
assign addr[43757]= 734482665;
assign addr[43758]= 805879757;
assign addr[43759]= 876254528;
assign addr[43760]= 945517704;
assign addr[43761]= 1013581418;
assign addr[43762]= 1080359326;
assign addr[43763]= 1145766716;
assign addr[43764]= 1209720613;
assign addr[43765]= 1272139887;
assign addr[43766]= 1332945355;
assign addr[43767]= 1392059879;
assign addr[43768]= 1449408469;
assign addr[43769]= 1504918373;
assign addr[43770]= 1558519173;
assign addr[43771]= 1610142873;
assign addr[43772]= 1659723983;
assign addr[43773]= 1707199606;
assign addr[43774]= 1752509516;
assign addr[43775]= 1795596234;
assign addr[43776]= 1836405100;
assign addr[43777]= 1874884346;
assign addr[43778]= 1910985158;
assign addr[43779]= 1944661739;
assign addr[43780]= 1975871368;
assign addr[43781]= 2004574453;
assign addr[43782]= 2030734582;
assign addr[43783]= 2054318569;
assign addr[43784]= 2075296495;
assign addr[43785]= 2093641749;
assign addr[43786]= 2109331059;
assign addr[43787]= 2122344521;
assign addr[43788]= 2132665626;
assign addr[43789]= 2140281282;
assign addr[43790]= 2145181827;
assign addr[43791]= 2147361045;
assign addr[43792]= 2146816171;
assign addr[43793]= 2143547897;
assign addr[43794]= 2137560369;
assign addr[43795]= 2128861181;
assign addr[43796]= 2117461370;
assign addr[43797]= 2103375398;
assign addr[43798]= 2086621133;
assign addr[43799]= 2067219829;
assign addr[43800]= 2045196100;
assign addr[43801]= 2020577882;
assign addr[43802]= 1993396407;
assign addr[43803]= 1963686155;
assign addr[43804]= 1931484818;
assign addr[43805]= 1896833245;
assign addr[43806]= 1859775393;
assign addr[43807]= 1820358275;
assign addr[43808]= 1778631892;
assign addr[43809]= 1734649179;
assign addr[43810]= 1688465931;
assign addr[43811]= 1640140734;
assign addr[43812]= 1589734894;
assign addr[43813]= 1537312353;
assign addr[43814]= 1482939614;
assign addr[43815]= 1426685652;
assign addr[43816]= 1368621831;
assign addr[43817]= 1308821808;
assign addr[43818]= 1247361445;
assign addr[43819]= 1184318708;
assign addr[43820]= 1119773573;
assign addr[43821]= 1053807919;
assign addr[43822]= 986505429;
assign addr[43823]= 917951481;
assign addr[43824]= 848233042;
assign addr[43825]= 777438554;
assign addr[43826]= 705657826;
assign addr[43827]= 632981917;
assign addr[43828]= 559503022;
assign addr[43829]= 485314355;
assign addr[43830]= 410510029;
assign addr[43831]= 335184940;
assign addr[43832]= 259434643;
assign addr[43833]= 183355234;
assign addr[43834]= 107043224;
assign addr[43835]= 30595422;
assign addr[43836]= -45891193;
assign addr[43837]= -122319591;
assign addr[43838]= -198592817;
assign addr[43839]= -274614114;
assign addr[43840]= -350287041;
assign addr[43841]= -425515602;
assign addr[43842]= -500204365;
assign addr[43843]= -574258580;
assign addr[43844]= -647584304;
assign addr[43845]= -720088517;
assign addr[43846]= -791679244;
assign addr[43847]= -862265664;
assign addr[43848]= -931758235;
assign addr[43849]= -1000068799;
assign addr[43850]= -1067110699;
assign addr[43851]= -1132798888;
assign addr[43852]= -1197050035;
assign addr[43853]= -1259782632;
assign addr[43854]= -1320917099;
assign addr[43855]= -1380375881;
assign addr[43856]= -1438083551;
assign addr[43857]= -1493966902;
assign addr[43858]= -1547955041;
assign addr[43859]= -1599979481;
assign addr[43860]= -1649974225;
assign addr[43861]= -1697875851;
assign addr[43862]= -1743623590;
assign addr[43863]= -1787159411;
assign addr[43864]= -1828428082;
assign addr[43865]= -1867377253;
assign addr[43866]= -1903957513;
assign addr[43867]= -1938122457;
assign addr[43868]= -1969828744;
assign addr[43869]= -1999036154;
assign addr[43870]= -2025707632;
assign addr[43871]= -2049809346;
assign addr[43872]= -2071310720;
assign addr[43873]= -2090184478;
assign addr[43874]= -2106406677;
assign addr[43875]= -2119956737;
assign addr[43876]= -2130817471;
assign addr[43877]= -2138975100;
assign addr[43878]= -2144419275;
assign addr[43879]= -2147143090;
assign addr[43880]= -2147143090;
assign addr[43881]= -2144419275;
assign addr[43882]= -2138975100;
assign addr[43883]= -2130817471;
assign addr[43884]= -2119956737;
assign addr[43885]= -2106406677;
assign addr[43886]= -2090184478;
assign addr[43887]= -2071310720;
assign addr[43888]= -2049809346;
assign addr[43889]= -2025707632;
assign addr[43890]= -1999036154;
assign addr[43891]= -1969828744;
assign addr[43892]= -1938122457;
assign addr[43893]= -1903957513;
assign addr[43894]= -1867377253;
assign addr[43895]= -1828428082;
assign addr[43896]= -1787159411;
assign addr[43897]= -1743623590;
assign addr[43898]= -1697875851;
assign addr[43899]= -1649974225;
assign addr[43900]= -1599979481;
assign addr[43901]= -1547955041;
assign addr[43902]= -1493966902;
assign addr[43903]= -1438083551;
assign addr[43904]= -1380375881;
assign addr[43905]= -1320917099;
assign addr[43906]= -1259782632;
assign addr[43907]= -1197050035;
assign addr[43908]= -1132798888;
assign addr[43909]= -1067110699;
assign addr[43910]= -1000068799;
assign addr[43911]= -931758235;
assign addr[43912]= -862265664;
assign addr[43913]= -791679244;
assign addr[43914]= -720088517;
assign addr[43915]= -647584304;
assign addr[43916]= -574258580;
assign addr[43917]= -500204365;
assign addr[43918]= -425515602;
assign addr[43919]= -350287041;
assign addr[43920]= -274614114;
assign addr[43921]= -198592817;
assign addr[43922]= -122319591;
assign addr[43923]= -45891193;
assign addr[43924]= 30595422;
assign addr[43925]= 107043224;
assign addr[43926]= 183355234;
assign addr[43927]= 259434643;
assign addr[43928]= 335184940;
assign addr[43929]= 410510029;
assign addr[43930]= 485314355;
assign addr[43931]= 559503022;
assign addr[43932]= 632981917;
assign addr[43933]= 705657826;
assign addr[43934]= 777438554;
assign addr[43935]= 848233042;
assign addr[43936]= 917951481;
assign addr[43937]= 986505429;
assign addr[43938]= 1053807919;
assign addr[43939]= 1119773573;
assign addr[43940]= 1184318708;
assign addr[43941]= 1247361445;
assign addr[43942]= 1308821808;
assign addr[43943]= 1368621831;
assign addr[43944]= 1426685652;
assign addr[43945]= 1482939614;
assign addr[43946]= 1537312353;
assign addr[43947]= 1589734894;
assign addr[43948]= 1640140734;
assign addr[43949]= 1688465931;
assign addr[43950]= 1734649179;
assign addr[43951]= 1778631892;
assign addr[43952]= 1820358275;
assign addr[43953]= 1859775393;
assign addr[43954]= 1896833245;
assign addr[43955]= 1931484818;
assign addr[43956]= 1963686155;
assign addr[43957]= 1993396407;
assign addr[43958]= 2020577882;
assign addr[43959]= 2045196100;
assign addr[43960]= 2067219829;
assign addr[43961]= 2086621133;
assign addr[43962]= 2103375398;
assign addr[43963]= 2117461370;
assign addr[43964]= 2128861181;
assign addr[43965]= 2137560369;
assign addr[43966]= 2143547897;
assign addr[43967]= 2146816171;
assign addr[43968]= 2147361045;
assign addr[43969]= 2145181827;
assign addr[43970]= 2140281282;
assign addr[43971]= 2132665626;
assign addr[43972]= 2122344521;
assign addr[43973]= 2109331059;
assign addr[43974]= 2093641749;
assign addr[43975]= 2075296495;
assign addr[43976]= 2054318569;
assign addr[43977]= 2030734582;
assign addr[43978]= 2004574453;
assign addr[43979]= 1975871368;
assign addr[43980]= 1944661739;
assign addr[43981]= 1910985158;
assign addr[43982]= 1874884346;
assign addr[43983]= 1836405100;
assign addr[43984]= 1795596234;
assign addr[43985]= 1752509516;
assign addr[43986]= 1707199606;
assign addr[43987]= 1659723983;
assign addr[43988]= 1610142873;
assign addr[43989]= 1558519173;
assign addr[43990]= 1504918373;
assign addr[43991]= 1449408469;
assign addr[43992]= 1392059879;
assign addr[43993]= 1332945355;
assign addr[43994]= 1272139887;
assign addr[43995]= 1209720613;
assign addr[43996]= 1145766716;
assign addr[43997]= 1080359326;
assign addr[43998]= 1013581418;
assign addr[43999]= 945517704;
assign addr[44000]= 876254528;
assign addr[44001]= 805879757;
assign addr[44002]= 734482665;
assign addr[44003]= 662153826;
assign addr[44004]= 588984994;
assign addr[44005]= 515068990;
assign addr[44006]= 440499581;
assign addr[44007]= 365371365;
assign addr[44008]= 289779648;
assign addr[44009]= 213820322;
assign addr[44010]= 137589750;
assign addr[44011]= 61184634;
assign addr[44012]= -15298099;
assign addr[44013]= -91761426;
assign addr[44014]= -168108346;
assign addr[44015]= -244242007;
assign addr[44016]= -320065829;
assign addr[44017]= -395483624;
assign addr[44018]= -470399716;
assign addr[44019]= -544719071;
assign addr[44020]= -618347408;
assign addr[44021]= -691191324;
assign addr[44022]= -763158411;
assign addr[44023]= -834157373;
assign addr[44024]= -904098143;
assign addr[44025]= -972891995;
assign addr[44026]= -1040451659;
assign addr[44027]= -1106691431;
assign addr[44028]= -1171527280;
assign addr[44029]= -1234876957;
assign addr[44030]= -1296660098;
assign addr[44031]= -1356798326;
assign addr[44032]= -1415215352;
assign addr[44033]= -1471837070;
assign addr[44034]= -1526591649;
assign addr[44035]= -1579409630;
assign addr[44036]= -1630224009;
assign addr[44037]= -1678970324;
assign addr[44038]= -1725586737;
assign addr[44039]= -1770014111;
assign addr[44040]= -1812196087;
assign addr[44041]= -1852079154;
assign addr[44042]= -1889612716;
assign addr[44043]= -1924749160;
assign addr[44044]= -1957443913;
assign addr[44045]= -1987655498;
assign addr[44046]= -2015345591;
assign addr[44047]= -2040479063;
assign addr[44048]= -2063024031;
assign addr[44049]= -2082951896;
assign addr[44050]= -2100237377;
assign addr[44051]= -2114858546;
assign addr[44052]= -2126796855;
assign addr[44053]= -2136037160;
assign addr[44054]= -2142567738;
assign addr[44055]= -2146380306;
assign addr[44056]= -2147470025;
assign addr[44057]= -2145835515;
assign addr[44058]= -2141478848;
assign addr[44059]= -2134405552;
assign addr[44060]= -2124624598;
assign addr[44061]= -2112148396;
assign addr[44062]= -2096992772;
assign addr[44063]= -2079176953;
assign addr[44064]= -2058723538;
assign addr[44065]= -2035658475;
assign addr[44066]= -2010011024;
assign addr[44067]= -1981813720;
assign addr[44068]= -1951102334;
assign addr[44069]= -1917915825;
assign addr[44070]= -1882296293;
assign addr[44071]= -1844288924;
assign addr[44072]= -1803941934;
assign addr[44073]= -1761306505;
assign addr[44074]= -1716436725;
assign addr[44075]= -1669389513;
assign addr[44076]= -1620224553;
assign addr[44077]= -1569004214;
assign addr[44078]= -1515793473;
assign addr[44079]= -1460659832;
assign addr[44080]= -1403673233;
assign addr[44081]= -1344905966;
assign addr[44082]= -1284432584;
assign addr[44083]= -1222329801;
assign addr[44084]= -1158676398;
assign addr[44085]= -1093553126;
assign addr[44086]= -1027042599;
assign addr[44087]= -959229189;
assign addr[44088]= -890198924;
assign addr[44089]= -820039373;
assign addr[44090]= -748839539;
assign addr[44091]= -676689746;
assign addr[44092]= -603681519;
assign addr[44093]= -529907477;
assign addr[44094]= -455461206;
assign addr[44095]= -380437148;
assign addr[44096]= -304930476;
assign addr[44097]= -229036977;
assign addr[44098]= -152852926;
assign addr[44099]= -76474970;
assign addr[44100]= 0;
assign addr[44101]= 76474970;
assign addr[44102]= 152852926;
assign addr[44103]= 229036977;
assign addr[44104]= 304930476;
assign addr[44105]= 380437148;
assign addr[44106]= 455461206;
assign addr[44107]= 529907477;
assign addr[44108]= 603681519;
assign addr[44109]= 676689746;
assign addr[44110]= 748839539;
assign addr[44111]= 820039373;
assign addr[44112]= 890198924;
assign addr[44113]= 959229189;
assign addr[44114]= 1027042599;
assign addr[44115]= 1093553126;
assign addr[44116]= 1158676398;
assign addr[44117]= 1222329801;
assign addr[44118]= 1284432584;
assign addr[44119]= 1344905966;
assign addr[44120]= 1403673233;
assign addr[44121]= 1460659832;
assign addr[44122]= 1515793473;
assign addr[44123]= 1569004214;
assign addr[44124]= 1620224553;
assign addr[44125]= 1669389513;
assign addr[44126]= 1716436725;
assign addr[44127]= 1761306505;
assign addr[44128]= 1803941934;
assign addr[44129]= 1844288924;
assign addr[44130]= 1882296293;
assign addr[44131]= 1917915825;
assign addr[44132]= 1951102334;
assign addr[44133]= 1981813720;
assign addr[44134]= 2010011024;
assign addr[44135]= 2035658475;
assign addr[44136]= 2058723538;
assign addr[44137]= 2079176953;
assign addr[44138]= 2096992772;
assign addr[44139]= 2112148396;
assign addr[44140]= 2124624598;
assign addr[44141]= 2134405552;
assign addr[44142]= 2141478848;
assign addr[44143]= 2145835515;
assign addr[44144]= 2147470025;
assign addr[44145]= 2146380306;
assign addr[44146]= 2142567738;
assign addr[44147]= 2136037160;
assign addr[44148]= 2126796855;
assign addr[44149]= 2114858546;
assign addr[44150]= 2100237377;
assign addr[44151]= 2082951896;
assign addr[44152]= 2063024031;
assign addr[44153]= 2040479063;
assign addr[44154]= 2015345591;
assign addr[44155]= 1987655498;
assign addr[44156]= 1957443913;
assign addr[44157]= 1924749160;
assign addr[44158]= 1889612716;
assign addr[44159]= 1852079154;
assign addr[44160]= 1812196087;
assign addr[44161]= 1770014111;
assign addr[44162]= 1725586737;
assign addr[44163]= 1678970324;
assign addr[44164]= 1630224009;
assign addr[44165]= 1579409630;
assign addr[44166]= 1526591649;
assign addr[44167]= 1471837070;
assign addr[44168]= 1415215352;
assign addr[44169]= 1356798326;
assign addr[44170]= 1296660098;
assign addr[44171]= 1234876957;
assign addr[44172]= 1171527280;
assign addr[44173]= 1106691431;
assign addr[44174]= 1040451659;
assign addr[44175]= 972891995;
assign addr[44176]= 904098143;
assign addr[44177]= 834157373;
assign addr[44178]= 763158411;
assign addr[44179]= 691191324;
assign addr[44180]= 618347408;
assign addr[44181]= 544719071;
assign addr[44182]= 470399716;
assign addr[44183]= 395483624;
assign addr[44184]= 320065829;
assign addr[44185]= 244242007;
assign addr[44186]= 168108346;
assign addr[44187]= 91761426;
assign addr[44188]= 15298099;
assign addr[44189]= -61184634;
assign addr[44190]= -137589750;
assign addr[44191]= -213820322;
assign addr[44192]= -289779648;
assign addr[44193]= -365371365;
assign addr[44194]= -440499581;
assign addr[44195]= -515068990;
assign addr[44196]= -588984994;
assign addr[44197]= -662153826;
assign addr[44198]= -734482665;
assign addr[44199]= -805879757;
assign addr[44200]= -876254528;
assign addr[44201]= -945517704;
assign addr[44202]= -1013581418;
assign addr[44203]= -1080359326;
assign addr[44204]= -1145766716;
assign addr[44205]= -1209720613;
assign addr[44206]= -1272139887;
assign addr[44207]= -1332945355;
assign addr[44208]= -1392059879;
assign addr[44209]= -1449408469;
assign addr[44210]= -1504918373;
assign addr[44211]= -1558519173;
assign addr[44212]= -1610142873;
assign addr[44213]= -1659723983;
assign addr[44214]= -1707199606;
assign addr[44215]= -1752509516;
assign addr[44216]= -1795596234;
assign addr[44217]= -1836405100;
assign addr[44218]= -1874884346;
assign addr[44219]= -1910985158;
assign addr[44220]= -1944661739;
assign addr[44221]= -1975871368;
assign addr[44222]= -2004574453;
assign addr[44223]= -2030734582;
assign addr[44224]= -2054318569;
assign addr[44225]= -2075296495;
assign addr[44226]= -2093641749;
assign addr[44227]= -2109331059;
assign addr[44228]= -2122344521;
assign addr[44229]= -2132665626;
assign addr[44230]= -2140281282;
assign addr[44231]= -2145181827;
assign addr[44232]= -2147361045;
assign addr[44233]= -2146816171;
assign addr[44234]= -2143547897;
assign addr[44235]= -2137560369;
assign addr[44236]= -2128861181;
assign addr[44237]= -2117461370;
assign addr[44238]= -2103375398;
assign addr[44239]= -2086621133;
assign addr[44240]= -2067219829;
assign addr[44241]= -2045196100;
assign addr[44242]= -2020577882;
assign addr[44243]= -1993396407;
assign addr[44244]= -1963686155;
assign addr[44245]= -1931484818;
assign addr[44246]= -1896833245;
assign addr[44247]= -1859775393;
assign addr[44248]= -1820358275;
assign addr[44249]= -1778631892;
assign addr[44250]= -1734649179;
assign addr[44251]= -1688465931;
assign addr[44252]= -1640140734;
assign addr[44253]= -1589734894;
assign addr[44254]= -1537312353;
assign addr[44255]= -1482939614;
assign addr[44256]= -1426685652;
assign addr[44257]= -1368621831;
assign addr[44258]= -1308821808;
assign addr[44259]= -1247361445;
assign addr[44260]= -1184318708;
assign addr[44261]= -1119773573;
assign addr[44262]= -1053807919;
assign addr[44263]= -986505429;
assign addr[44264]= -917951481;
assign addr[44265]= -848233042;
assign addr[44266]= -777438554;
assign addr[44267]= -705657826;
assign addr[44268]= -632981917;
assign addr[44269]= -559503022;
assign addr[44270]= -485314355;
assign addr[44271]= -410510029;
assign addr[44272]= -335184940;
assign addr[44273]= -259434643;
assign addr[44274]= -183355234;
assign addr[44275]= -107043224;
assign addr[44276]= -30595422;
assign addr[44277]= 45891193;
assign addr[44278]= 122319591;
assign addr[44279]= 198592817;
assign addr[44280]= 274614114;
assign addr[44281]= 350287041;
assign addr[44282]= 425515602;
assign addr[44283]= 500204365;
assign addr[44284]= 574258580;
assign addr[44285]= 647584304;
assign addr[44286]= 720088517;
assign addr[44287]= 791679244;
assign addr[44288]= 862265664;
assign addr[44289]= 931758235;
assign addr[44290]= 1000068799;
assign addr[44291]= 1067110699;
assign addr[44292]= 1132798888;
assign addr[44293]= 1197050035;
assign addr[44294]= 1259782632;
assign addr[44295]= 1320917099;
assign addr[44296]= 1380375881;
assign addr[44297]= 1438083551;
assign addr[44298]= 1493966902;
assign addr[44299]= 1547955041;
assign addr[44300]= 1599979481;
assign addr[44301]= 1649974225;
assign addr[44302]= 1697875851;
assign addr[44303]= 1743623590;
assign addr[44304]= 1787159411;
assign addr[44305]= 1828428082;
assign addr[44306]= 1867377253;
assign addr[44307]= 1903957513;
assign addr[44308]= 1938122457;
assign addr[44309]= 1969828744;
assign addr[44310]= 1999036154;
assign addr[44311]= 2025707632;
assign addr[44312]= 2049809346;
assign addr[44313]= 2071310720;
assign addr[44314]= 2090184478;
assign addr[44315]= 2106406677;
assign addr[44316]= 2119956737;
assign addr[44317]= 2130817471;
assign addr[44318]= 2138975100;
assign addr[44319]= 2144419275;
assign addr[44320]= 2147143090;
assign addr[44321]= 2147143090;
assign addr[44322]= 2144419275;
assign addr[44323]= 2138975100;
assign addr[44324]= 2130817471;
assign addr[44325]= 2119956737;
assign addr[44326]= 2106406677;
assign addr[44327]= 2090184478;
assign addr[44328]= 2071310720;
assign addr[44329]= 2049809346;
assign addr[44330]= 2025707632;
assign addr[44331]= 1999036154;
assign addr[44332]= 1969828744;
assign addr[44333]= 1938122457;
assign addr[44334]= 1903957513;
assign addr[44335]= 1867377253;
assign addr[44336]= 1828428082;
assign addr[44337]= 1787159411;
assign addr[44338]= 1743623590;
assign addr[44339]= 1697875851;
assign addr[44340]= 1649974225;
assign addr[44341]= 1599979481;
assign addr[44342]= 1547955041;
assign addr[44343]= 1493966902;
assign addr[44344]= 1438083551;
assign addr[44345]= 1380375881;
assign addr[44346]= 1320917099;
assign addr[44347]= 1259782632;
assign addr[44348]= 1197050035;
assign addr[44349]= 1132798888;
assign addr[44350]= 1067110699;
assign addr[44351]= 1000068799;
assign addr[44352]= 931758235;
assign addr[44353]= 862265664;
assign addr[44354]= 791679244;
assign addr[44355]= 720088517;
assign addr[44356]= 647584304;
assign addr[44357]= 574258580;
assign addr[44358]= 500204365;
assign addr[44359]= 425515602;
assign addr[44360]= 350287041;
assign addr[44361]= 274614114;
assign addr[44362]= 198592817;
assign addr[44363]= 122319591;
assign addr[44364]= 45891193;
assign addr[44365]= -30595422;
assign addr[44366]= -107043224;
assign addr[44367]= -183355234;
assign addr[44368]= -259434643;
assign addr[44369]= -335184940;
assign addr[44370]= -410510029;
assign addr[44371]= -485314355;
assign addr[44372]= -559503022;
assign addr[44373]= -632981917;
assign addr[44374]= -705657826;
assign addr[44375]= -777438554;
assign addr[44376]= -848233042;
assign addr[44377]= -917951481;
assign addr[44378]= -986505429;
assign addr[44379]= -1053807919;
assign addr[44380]= -1119773573;
assign addr[44381]= -1184318708;
assign addr[44382]= -1247361445;
assign addr[44383]= -1308821808;
assign addr[44384]= -1368621831;
assign addr[44385]= -1426685652;
assign addr[44386]= -1482939614;
assign addr[44387]= -1537312353;
assign addr[44388]= -1589734894;
assign addr[44389]= -1640140734;
assign addr[44390]= -1688465931;
assign addr[44391]= -1734649179;
assign addr[44392]= -1778631892;
assign addr[44393]= -1820358275;
assign addr[44394]= -1859775393;
assign addr[44395]= -1896833245;
assign addr[44396]= -1931484818;
assign addr[44397]= -1963686155;
assign addr[44398]= -1993396407;
assign addr[44399]= -2020577882;
assign addr[44400]= -2045196100;
assign addr[44401]= -2067219829;
assign addr[44402]= -2086621133;
assign addr[44403]= -2103375398;
assign addr[44404]= -2117461370;
assign addr[44405]= -2128861181;
assign addr[44406]= -2137560369;
assign addr[44407]= -2143547897;
assign addr[44408]= -2146816171;
assign addr[44409]= -2147361045;
assign addr[44410]= -2145181827;
assign addr[44411]= -2140281282;
assign addr[44412]= -2132665626;
assign addr[44413]= -2122344521;
assign addr[44414]= -2109331059;
assign addr[44415]= -2093641749;
assign addr[44416]= -2075296495;
assign addr[44417]= -2054318569;
assign addr[44418]= -2030734582;
assign addr[44419]= -2004574453;
assign addr[44420]= -1975871368;
assign addr[44421]= -1944661739;
assign addr[44422]= -1910985158;
assign addr[44423]= -1874884346;
assign addr[44424]= -1836405100;
assign addr[44425]= -1795596234;
assign addr[44426]= -1752509516;
assign addr[44427]= -1707199606;
assign addr[44428]= -1659723983;
assign addr[44429]= -1610142873;
assign addr[44430]= -1558519173;
assign addr[44431]= -1504918373;
assign addr[44432]= -1449408469;
assign addr[44433]= -1392059879;
assign addr[44434]= -1332945355;
assign addr[44435]= -1272139887;
assign addr[44436]= -1209720613;
assign addr[44437]= -1145766716;
assign addr[44438]= -1080359326;
assign addr[44439]= -1013581418;
assign addr[44440]= -945517704;
assign addr[44441]= -876254528;
assign addr[44442]= -805879757;
assign addr[44443]= -734482665;
assign addr[44444]= -662153826;
assign addr[44445]= -588984994;
assign addr[44446]= -515068990;
assign addr[44447]= -440499581;
assign addr[44448]= -365371365;
assign addr[44449]= -289779648;
assign addr[44450]= -213820322;
assign addr[44451]= -137589750;
assign addr[44452]= -61184634;
assign addr[44453]= 15298099;
assign addr[44454]= 91761426;
assign addr[44455]= 168108346;
assign addr[44456]= 244242007;
assign addr[44457]= 320065829;
assign addr[44458]= 395483624;
assign addr[44459]= 470399716;
assign addr[44460]= 544719071;
assign addr[44461]= 618347408;
assign addr[44462]= 691191324;
assign addr[44463]= 763158411;
assign addr[44464]= 834157373;
assign addr[44465]= 904098143;
assign addr[44466]= 972891995;
assign addr[44467]= 1040451659;
assign addr[44468]= 1106691431;
assign addr[44469]= 1171527280;
assign addr[44470]= 1234876957;
assign addr[44471]= 1296660098;
assign addr[44472]= 1356798326;
assign addr[44473]= 1415215352;
assign addr[44474]= 1471837070;
assign addr[44475]= 1526591649;
assign addr[44476]= 1579409630;
assign addr[44477]= 1630224009;
assign addr[44478]= 1678970324;
assign addr[44479]= 1725586737;
assign addr[44480]= 1770014111;
assign addr[44481]= 1812196087;
assign addr[44482]= 1852079154;
assign addr[44483]= 1889612716;
assign addr[44484]= 1924749160;
assign addr[44485]= 1957443913;
assign addr[44486]= 1987655498;
assign addr[44487]= 2015345591;
assign addr[44488]= 2040479063;
assign addr[44489]= 2063024031;
assign addr[44490]= 2082951896;
assign addr[44491]= 2100237377;
assign addr[44492]= 2114858546;
assign addr[44493]= 2126796855;
assign addr[44494]= 2136037160;
assign addr[44495]= 2142567738;
assign addr[44496]= 2146380306;
assign addr[44497]= 2147470025;
assign addr[44498]= 2145835515;
assign addr[44499]= 2141478848;
assign addr[44500]= 2134405552;
assign addr[44501]= 2124624598;
assign addr[44502]= 2112148396;
assign addr[44503]= 2096992772;
assign addr[44504]= 2079176953;
assign addr[44505]= 2058723538;
assign addr[44506]= 2035658475;
assign addr[44507]= 2010011024;
assign addr[44508]= 1981813720;
assign addr[44509]= 1951102334;
assign addr[44510]= 1917915825;
assign addr[44511]= 1882296293;
assign addr[44512]= 1844288924;
assign addr[44513]= 1803941934;
assign addr[44514]= 1761306505;
assign addr[44515]= 1716436725;
assign addr[44516]= 1669389513;
assign addr[44517]= 1620224553;
assign addr[44518]= 1569004214;
assign addr[44519]= 1515793473;
assign addr[44520]= 1460659832;
assign addr[44521]= 1403673233;
assign addr[44522]= 1344905966;
assign addr[44523]= 1284432584;
assign addr[44524]= 1222329801;
assign addr[44525]= 1158676398;
assign addr[44526]= 1093553126;
assign addr[44527]= 1027042599;
assign addr[44528]= 959229189;
assign addr[44529]= 890198924;
assign addr[44530]= 820039373;
assign addr[44531]= 748839539;
assign addr[44532]= 676689746;
assign addr[44533]= 603681519;
assign addr[44534]= 529907477;
assign addr[44535]= 455461206;
assign addr[44536]= 380437148;
assign addr[44537]= 304930476;
assign addr[44538]= 229036977;
assign addr[44539]= 152852926;
assign addr[44540]= 76474970;
assign addr[44541]= 0;
assign addr[44542]= -76474970;
assign addr[44543]= -152852926;
assign addr[44544]= -229036977;
assign addr[44545]= -304930476;
assign addr[44546]= -380437148;
assign addr[44547]= -455461206;
assign addr[44548]= -529907477;
assign addr[44549]= -603681519;
assign addr[44550]= -676689746;
assign addr[44551]= -748839539;
assign addr[44552]= -820039373;
assign addr[44553]= -890198924;
assign addr[44554]= -959229189;
assign addr[44555]= -1027042599;
assign addr[44556]= -1093553126;
assign addr[44557]= -1158676398;
assign addr[44558]= -1222329801;
assign addr[44559]= -1284432584;
assign addr[44560]= -1344905966;
assign addr[44561]= -1403673233;
assign addr[44562]= -1460659832;
assign addr[44563]= -1515793473;
assign addr[44564]= -1569004214;
assign addr[44565]= -1620224553;
assign addr[44566]= -1669389513;
assign addr[44567]= -1716436725;
assign addr[44568]= -1761306505;
assign addr[44569]= -1803941934;
assign addr[44570]= -1844288924;
assign addr[44571]= -1882296293;
assign addr[44572]= -1917915825;
assign addr[44573]= -1951102334;
assign addr[44574]= -1981813720;
assign addr[44575]= -2010011024;
assign addr[44576]= -2035658475;
assign addr[44577]= -2058723538;
assign addr[44578]= -2079176953;
assign addr[44579]= -2096992772;
assign addr[44580]= -2112148396;
assign addr[44581]= -2124624598;
assign addr[44582]= -2134405552;
assign addr[44583]= -2141478848;
assign addr[44584]= -2145835515;
assign addr[44585]= -2147470025;
assign addr[44586]= -2146380306;
assign addr[44587]= -2142567738;
assign addr[44588]= -2136037160;
assign addr[44589]= -2126796855;
assign addr[44590]= -2114858546;
assign addr[44591]= -2100237377;
assign addr[44592]= -2082951896;
assign addr[44593]= -2063024031;
assign addr[44594]= -2040479063;
assign addr[44595]= -2015345591;
assign addr[44596]= -1987655498;
assign addr[44597]= -1957443913;
assign addr[44598]= -1924749160;
assign addr[44599]= -1889612716;
assign addr[44600]= -1852079154;
assign addr[44601]= -1812196087;
assign addr[44602]= -1770014111;
assign addr[44603]= -1725586737;
assign addr[44604]= -1678970324;
assign addr[44605]= -1630224009;
assign addr[44606]= -1579409630;
assign addr[44607]= -1526591649;
assign addr[44608]= -1471837070;
assign addr[44609]= -1415215352;
assign addr[44610]= -1356798326;
assign addr[44611]= -1296660098;
assign addr[44612]= -1234876957;
assign addr[44613]= -1171527280;
assign addr[44614]= -1106691431;
assign addr[44615]= -1040451659;
assign addr[44616]= -972891995;
assign addr[44617]= -904098143;
assign addr[44618]= -834157373;
assign addr[44619]= -763158411;
assign addr[44620]= -691191324;
assign addr[44621]= -618347408;
assign addr[44622]= -544719071;
assign addr[44623]= -470399716;
assign addr[44624]= -395483624;
assign addr[44625]= -320065829;
assign addr[44626]= -244242007;
assign addr[44627]= -168108346;
assign addr[44628]= -91761426;
assign addr[44629]= -15298099;
assign addr[44630]= 61184634;
assign addr[44631]= 137589750;
assign addr[44632]= 213820322;
assign addr[44633]= 289779648;
assign addr[44634]= 365371365;
assign addr[44635]= 440499581;
assign addr[44636]= 515068990;
assign addr[44637]= 588984994;
assign addr[44638]= 662153826;
assign addr[44639]= 734482665;
assign addr[44640]= 805879757;
assign addr[44641]= 876254528;
assign addr[44642]= 945517704;
assign addr[44643]= 1013581418;
assign addr[44644]= 1080359326;
assign addr[44645]= 1145766716;
assign addr[44646]= 1209720613;
assign addr[44647]= 1272139887;
assign addr[44648]= 1332945355;
assign addr[44649]= 1392059879;
assign addr[44650]= 1449408469;
assign addr[44651]= 1504918373;
assign addr[44652]= 1558519173;
assign addr[44653]= 1610142873;
assign addr[44654]= 1659723983;
assign addr[44655]= 1707199606;
assign addr[44656]= 1752509516;
assign addr[44657]= 1795596234;
assign addr[44658]= 1836405100;
assign addr[44659]= 1874884346;
assign addr[44660]= 1910985158;
assign addr[44661]= 1944661739;
assign addr[44662]= 1975871368;
assign addr[44663]= 2004574453;
assign addr[44664]= 2030734582;
assign addr[44665]= 2054318569;
assign addr[44666]= 2075296495;
assign addr[44667]= 2093641749;
assign addr[44668]= 2109331059;
assign addr[44669]= 2122344521;
assign addr[44670]= 2132665626;
assign addr[44671]= 2140281282;
assign addr[44672]= 2145181827;
assign addr[44673]= 2147361045;
assign addr[44674]= 2146816171;
assign addr[44675]= 2143547897;
assign addr[44676]= 2137560369;
assign addr[44677]= 2128861181;
assign addr[44678]= 2117461370;
assign addr[44679]= 2103375398;
assign addr[44680]= 2086621133;
assign addr[44681]= 2067219829;
assign addr[44682]= 2045196100;
assign addr[44683]= 2020577882;
assign addr[44684]= 1993396407;
assign addr[44685]= 1963686155;
assign addr[44686]= 1931484818;
assign addr[44687]= 1896833245;
assign addr[44688]= 1859775393;
assign addr[44689]= 1820358275;
assign addr[44690]= 1778631892;
assign addr[44691]= 1734649179;
assign addr[44692]= 1688465931;
assign addr[44693]= 1640140734;
assign addr[44694]= 1589734894;
assign addr[44695]= 1537312353;
assign addr[44696]= 1482939614;
assign addr[44697]= 1426685652;
assign addr[44698]= 1368621831;
assign addr[44699]= 1308821808;
assign addr[44700]= 1247361445;
assign addr[44701]= 1184318708;
assign addr[44702]= 1119773573;
assign addr[44703]= 1053807919;
assign addr[44704]= 986505429;
assign addr[44705]= 917951481;
assign addr[44706]= 848233042;
assign addr[44707]= 777438554;
assign addr[44708]= 705657826;
assign addr[44709]= 632981917;
assign addr[44710]= 559503022;
assign addr[44711]= 485314355;
assign addr[44712]= 410510029;
assign addr[44713]= 335184940;
assign addr[44714]= 259434643;
assign addr[44715]= 183355234;
assign addr[44716]= 107043224;
assign addr[44717]= 30595422;
assign addr[44718]= -45891193;
assign addr[44719]= -122319591;
assign addr[44720]= -198592817;
assign addr[44721]= -274614114;
assign addr[44722]= -350287041;
assign addr[44723]= -425515602;
assign addr[44724]= -500204365;
assign addr[44725]= -574258580;
assign addr[44726]= -647584304;
assign addr[44727]= -720088517;
assign addr[44728]= -791679244;
assign addr[44729]= -862265664;
assign addr[44730]= -931758235;
assign addr[44731]= -1000068799;
assign addr[44732]= -1067110699;
assign addr[44733]= -1132798888;
assign addr[44734]= -1197050035;
assign addr[44735]= -1259782632;
assign addr[44736]= -1320917099;
assign addr[44737]= -1380375881;
assign addr[44738]= -1438083551;
assign addr[44739]= -1493966902;
assign addr[44740]= -1547955041;
assign addr[44741]= -1599979481;
assign addr[44742]= -1649974225;
assign addr[44743]= -1697875851;
assign addr[44744]= -1743623590;
assign addr[44745]= -1787159411;
assign addr[44746]= -1828428082;
assign addr[44747]= -1867377253;
assign addr[44748]= -1903957513;
assign addr[44749]= -1938122457;
assign addr[44750]= -1969828744;
assign addr[44751]= -1999036154;
assign addr[44752]= -2025707632;
assign addr[44753]= -2049809346;
assign addr[44754]= -2071310720;
assign addr[44755]= -2090184478;
assign addr[44756]= -2106406677;
assign addr[44757]= -2119956737;
assign addr[44758]= -2130817471;
assign addr[44759]= -2138975100;
assign addr[44760]= -2144419275;
assign addr[44761]= -2147143090;
assign addr[44762]= -2147143090;
assign addr[44763]= -2144419275;
assign addr[44764]= -2138975100;
assign addr[44765]= -2130817471;
assign addr[44766]= -2119956737;
assign addr[44767]= -2106406677;
assign addr[44768]= -2090184478;
assign addr[44769]= -2071310720;
assign addr[44770]= -2049809346;
assign addr[44771]= -2025707632;
assign addr[44772]= -1999036154;
assign addr[44773]= -1969828744;
assign addr[44774]= -1938122457;
assign addr[44775]= -1903957513;
assign addr[44776]= -1867377253;
assign addr[44777]= -1828428082;
assign addr[44778]= -1787159411;
assign addr[44779]= -1743623590;
assign addr[44780]= -1697875851;
assign addr[44781]= -1649974225;
assign addr[44782]= -1599979481;
assign addr[44783]= -1547955041;
assign addr[44784]= -1493966902;
assign addr[44785]= -1438083551;
assign addr[44786]= -1380375881;
assign addr[44787]= -1320917099;
assign addr[44788]= -1259782632;
assign addr[44789]= -1197050035;
assign addr[44790]= -1132798888;
assign addr[44791]= -1067110699;
assign addr[44792]= -1000068799;
assign addr[44793]= -931758235;
assign addr[44794]= -862265664;
assign addr[44795]= -791679244;
assign addr[44796]= -720088517;
assign addr[44797]= -647584304;
assign addr[44798]= -574258580;
assign addr[44799]= -500204365;
assign addr[44800]= -425515602;
assign addr[44801]= -350287041;
assign addr[44802]= -274614114;
assign addr[44803]= -198592817;
assign addr[44804]= -122319591;
assign addr[44805]= -45891193;
assign addr[44806]= 30595422;
assign addr[44807]= 107043224;
assign addr[44808]= 183355234;
assign addr[44809]= 259434643;
assign addr[44810]= 335184940;
assign addr[44811]= 410510029;
assign addr[44812]= 485314355;
assign addr[44813]= 559503022;
assign addr[44814]= 632981917;
assign addr[44815]= 705657826;
assign addr[44816]= 777438554;
assign addr[44817]= 848233042;
assign addr[44818]= 917951481;
assign addr[44819]= 986505429;
assign addr[44820]= 1053807919;
assign addr[44821]= 1119773573;
assign addr[44822]= 1184318708;
assign addr[44823]= 1247361445;
assign addr[44824]= 1308821808;
assign addr[44825]= 1368621831;
assign addr[44826]= 1426685652;
assign addr[44827]= 1482939614;
assign addr[44828]= 1537312353;
assign addr[44829]= 1589734894;
assign addr[44830]= 1640140734;
assign addr[44831]= 1688465931;
assign addr[44832]= 1734649179;
assign addr[44833]= 1778631892;
assign addr[44834]= 1820358275;
assign addr[44835]= 1859775393;
assign addr[44836]= 1896833245;
assign addr[44837]= 1931484818;
assign addr[44838]= 1963686155;
assign addr[44839]= 1993396407;
assign addr[44840]= 2020577882;
assign addr[44841]= 2045196100;
assign addr[44842]= 2067219829;
assign addr[44843]= 2086621133;
assign addr[44844]= 2103375398;
assign addr[44845]= 2117461370;
assign addr[44846]= 2128861181;
assign addr[44847]= 2137560369;
assign addr[44848]= 2143547897;
assign addr[44849]= 2146816171;
assign addr[44850]= 2147361045;
assign addr[44851]= 2145181827;
assign addr[44852]= 2140281282;
assign addr[44853]= 2132665626;
assign addr[44854]= 2122344521;
assign addr[44855]= 2109331059;
assign addr[44856]= 2093641749;
assign addr[44857]= 2075296495;
assign addr[44858]= 2054318569;
assign addr[44859]= 2030734582;
assign addr[44860]= 2004574453;
assign addr[44861]= 1975871368;
assign addr[44862]= 1944661739;
assign addr[44863]= 1910985158;
assign addr[44864]= 1874884346;
assign addr[44865]= 1836405100;
assign addr[44866]= 1795596234;
assign addr[44867]= 1752509516;
assign addr[44868]= 1707199606;
assign addr[44869]= 1659723983;
assign addr[44870]= 1610142873;
assign addr[44871]= 1558519173;
assign addr[44872]= 1504918373;
assign addr[44873]= 1449408469;
assign addr[44874]= 1392059879;
assign addr[44875]= 1332945355;
assign addr[44876]= 1272139887;
assign addr[44877]= 1209720613;
assign addr[44878]= 1145766716;
assign addr[44879]= 1080359326;
assign addr[44880]= 1013581418;
assign addr[44881]= 945517704;
assign addr[44882]= 876254528;
assign addr[44883]= 805879757;
assign addr[44884]= 734482665;
assign addr[44885]= 662153826;
assign addr[44886]= 588984994;
assign addr[44887]= 515068990;
assign addr[44888]= 440499581;
assign addr[44889]= 365371365;
assign addr[44890]= 289779648;
assign addr[44891]= 213820322;
assign addr[44892]= 137589750;
assign addr[44893]= 61184634;
assign addr[44894]= -15298099;
assign addr[44895]= -91761426;
assign addr[44896]= -168108346;
assign addr[44897]= -244242007;
assign addr[44898]= -320065829;
assign addr[44899]= -395483624;
assign addr[44900]= -470399716;
assign addr[44901]= -544719071;
assign addr[44902]= -618347408;
assign addr[44903]= -691191324;
assign addr[44904]= -763158411;
assign addr[44905]= -834157373;
assign addr[44906]= -904098143;
assign addr[44907]= -972891995;
assign addr[44908]= -1040451659;
assign addr[44909]= -1106691431;
assign addr[44910]= -1171527280;
assign addr[44911]= -1234876957;
assign addr[44912]= -1296660098;
assign addr[44913]= -1356798326;
assign addr[44914]= -1415215352;
assign addr[44915]= -1471837070;
assign addr[44916]= -1526591649;
assign addr[44917]= -1579409630;
assign addr[44918]= -1630224009;
assign addr[44919]= -1678970324;
assign addr[44920]= -1725586737;
assign addr[44921]= -1770014111;
assign addr[44922]= -1812196087;
assign addr[44923]= -1852079154;
assign addr[44924]= -1889612716;
assign addr[44925]= -1924749160;
assign addr[44926]= -1957443913;
assign addr[44927]= -1987655498;
assign addr[44928]= -2015345591;
assign addr[44929]= -2040479063;
assign addr[44930]= -2063024031;
assign addr[44931]= -2082951896;
assign addr[44932]= -2100237377;
assign addr[44933]= -2114858546;
assign addr[44934]= -2126796855;
assign addr[44935]= -2136037160;
assign addr[44936]= -2142567738;
assign addr[44937]= -2146380306;
assign addr[44938]= -2147470025;
assign addr[44939]= -2145835515;
assign addr[44940]= -2141478848;
assign addr[44941]= -2134405552;
assign addr[44942]= -2124624598;
assign addr[44943]= -2112148396;
assign addr[44944]= -2096992772;
assign addr[44945]= -2079176953;
assign addr[44946]= -2058723538;
assign addr[44947]= -2035658475;
assign addr[44948]= -2010011024;
assign addr[44949]= -1981813720;
assign addr[44950]= -1951102334;
assign addr[44951]= -1917915825;
assign addr[44952]= -1882296293;
assign addr[44953]= -1844288924;
assign addr[44954]= -1803941934;
assign addr[44955]= -1761306505;
assign addr[44956]= -1716436725;
assign addr[44957]= -1669389513;
assign addr[44958]= -1620224553;
assign addr[44959]= -1569004214;
assign addr[44960]= -1515793473;
assign addr[44961]= -1460659832;
assign addr[44962]= -1403673233;
assign addr[44963]= -1344905966;
assign addr[44964]= -1284432584;
assign addr[44965]= -1222329801;
assign addr[44966]= -1158676398;
assign addr[44967]= -1093553126;
assign addr[44968]= -1027042599;
assign addr[44969]= -959229189;
assign addr[44970]= -890198924;
assign addr[44971]= -820039373;
assign addr[44972]= -748839539;
assign addr[44973]= -676689746;
assign addr[44974]= -603681519;
assign addr[44975]= -529907477;
assign addr[44976]= -455461206;
assign addr[44977]= -380437148;
assign addr[44978]= -304930476;
assign addr[44979]= -229036977;
assign addr[44980]= -152852926;
assign addr[44981]= -76474970;
assign addr[44982]= 0;
assign addr[44983]= 76474970;
assign addr[44984]= 152852926;
assign addr[44985]= 229036977;
assign addr[44986]= 304930476;
assign addr[44987]= 380437148;
assign addr[44988]= 455461206;
assign addr[44989]= 529907477;
assign addr[44990]= 603681519;
assign addr[44991]= 676689746;
assign addr[44992]= 748839539;
assign addr[44993]= 820039373;
assign addr[44994]= 890198924;
assign addr[44995]= 959229189;
assign addr[44996]= 1027042599;
assign addr[44997]= 1093553126;
assign addr[44998]= 1158676398;
assign addr[44999]= 1222329801;
assign addr[45000]= 1284432584;
assign addr[45001]= 1344905966;
assign addr[45002]= 1403673233;
assign addr[45003]= 1460659832;
assign addr[45004]= 1515793473;
assign addr[45005]= 1569004214;
assign addr[45006]= 1620224553;
assign addr[45007]= 1669389513;
assign addr[45008]= 1716436725;
assign addr[45009]= 1761306505;
assign addr[45010]= 1803941934;
assign addr[45011]= 1844288924;
assign addr[45012]= 1882296293;
assign addr[45013]= 1917915825;
assign addr[45014]= 1951102334;
assign addr[45015]= 1981813720;
assign addr[45016]= 2010011024;
assign addr[45017]= 2035658475;
assign addr[45018]= 2058723538;
assign addr[45019]= 2079176953;
assign addr[45020]= 2096992772;
assign addr[45021]= 2112148396;
assign addr[45022]= 2124624598;
assign addr[45023]= 2134405552;
assign addr[45024]= 2141478848;
assign addr[45025]= 2145835515;
assign addr[45026]= 2147470025;
assign addr[45027]= 2146380306;
assign addr[45028]= 2142567738;
assign addr[45029]= 2136037160;
assign addr[45030]= 2126796855;
assign addr[45031]= 2114858546;
assign addr[45032]= 2100237377;
assign addr[45033]= 2082951896;
assign addr[45034]= 2063024031;
assign addr[45035]= 2040479063;
assign addr[45036]= 2015345591;
assign addr[45037]= 1987655498;
assign addr[45038]= 1957443913;
assign addr[45039]= 1924749160;
assign addr[45040]= 1889612716;
assign addr[45041]= 1852079154;
assign addr[45042]= 1812196087;
assign addr[45043]= 1770014111;
assign addr[45044]= 1725586737;
assign addr[45045]= 1678970324;
assign addr[45046]= 1630224009;
assign addr[45047]= 1579409630;
assign addr[45048]= 1526591649;
assign addr[45049]= 1471837070;
assign addr[45050]= 1415215352;
assign addr[45051]= 1356798326;
assign addr[45052]= 1296660098;
assign addr[45053]= 1234876957;
assign addr[45054]= 1171527280;
assign addr[45055]= 1106691431;
assign addr[45056]= 1040451659;
assign addr[45057]= 972891995;
assign addr[45058]= 904098143;
assign addr[45059]= 834157373;
assign addr[45060]= 763158411;
assign addr[45061]= 691191324;
assign addr[45062]= 618347408;
assign addr[45063]= 544719071;
assign addr[45064]= 470399716;
assign addr[45065]= 395483624;
assign addr[45066]= 320065829;
assign addr[45067]= 244242007;
assign addr[45068]= 168108346;
assign addr[45069]= 91761426;
assign addr[45070]= 15298099;
assign addr[45071]= -61184634;
assign addr[45072]= -137589750;
assign addr[45073]= -213820322;
assign addr[45074]= -289779648;
assign addr[45075]= -365371365;
assign addr[45076]= -440499581;
assign addr[45077]= -515068990;
assign addr[45078]= -588984994;
assign addr[45079]= -662153826;
assign addr[45080]= -734482665;
assign addr[45081]= -805879757;
assign addr[45082]= -876254528;
assign addr[45083]= -945517704;
assign addr[45084]= -1013581418;
assign addr[45085]= -1080359326;
assign addr[45086]= -1145766716;
assign addr[45087]= -1209720613;
assign addr[45088]= -1272139887;
assign addr[45089]= -1332945355;
assign addr[45090]= -1392059879;
assign addr[45091]= -1449408469;
assign addr[45092]= -1504918373;
assign addr[45093]= -1558519173;
assign addr[45094]= -1610142873;
assign addr[45095]= -1659723983;
assign addr[45096]= -1707199606;
assign addr[45097]= -1752509516;
assign addr[45098]= -1795596234;
assign addr[45099]= -1836405100;
assign addr[45100]= -1874884346;
assign addr[45101]= -1910985158;
assign addr[45102]= -1944661739;
assign addr[45103]= -1975871368;
assign addr[45104]= -2004574453;
assign addr[45105]= -2030734582;
assign addr[45106]= -2054318569;
assign addr[45107]= -2075296495;
assign addr[45108]= -2093641749;
assign addr[45109]= -2109331059;
assign addr[45110]= -2122344521;
assign addr[45111]= -2132665626;
assign addr[45112]= -2140281282;
assign addr[45113]= -2145181827;
assign addr[45114]= -2147361045;
assign addr[45115]= -2146816171;
assign addr[45116]= -2143547897;
assign addr[45117]= -2137560369;
assign addr[45118]= -2128861181;
assign addr[45119]= -2117461370;
assign addr[45120]= -2103375398;
assign addr[45121]= -2086621133;
assign addr[45122]= -2067219829;
assign addr[45123]= -2045196100;
assign addr[45124]= -2020577882;
assign addr[45125]= -1993396407;
assign addr[45126]= -1963686155;
assign addr[45127]= -1931484818;
assign addr[45128]= -1896833245;
assign addr[45129]= -1859775393;
assign addr[45130]= -1820358275;
assign addr[45131]= -1778631892;
assign addr[45132]= -1734649179;
assign addr[45133]= -1688465931;
assign addr[45134]= -1640140734;
assign addr[45135]= -1589734894;
assign addr[45136]= -1537312353;
assign addr[45137]= -1482939614;
assign addr[45138]= -1426685652;
assign addr[45139]= -1368621831;
assign addr[45140]= -1308821808;
assign addr[45141]= -1247361445;
assign addr[45142]= -1184318708;
assign addr[45143]= -1119773573;
assign addr[45144]= -1053807919;
assign addr[45145]= -986505429;
assign addr[45146]= -917951481;
assign addr[45147]= -848233042;
assign addr[45148]= -777438554;
assign addr[45149]= -705657826;
assign addr[45150]= -632981917;
assign addr[45151]= -559503022;
assign addr[45152]= -485314355;
assign addr[45153]= -410510029;
assign addr[45154]= -335184940;
assign addr[45155]= -259434643;
assign addr[45156]= -183355234;
assign addr[45157]= -107043224;
assign addr[45158]= -30595422;
assign addr[45159]= 45891193;
assign addr[45160]= 122319591;
assign addr[45161]= 198592817;
assign addr[45162]= 274614114;
assign addr[45163]= 350287041;
assign addr[45164]= 425515602;
assign addr[45165]= 500204365;
assign addr[45166]= 574258580;
assign addr[45167]= 647584304;
assign addr[45168]= 720088517;
assign addr[45169]= 791679244;
assign addr[45170]= 862265664;
assign addr[45171]= 931758235;
assign addr[45172]= 1000068799;
assign addr[45173]= 1067110699;
assign addr[45174]= 1132798888;
assign addr[45175]= 1197050035;
assign addr[45176]= 1259782632;
assign addr[45177]= 1320917099;
assign addr[45178]= 1380375881;
assign addr[45179]= 1438083551;
assign addr[45180]= 1493966902;
assign addr[45181]= 1547955041;
assign addr[45182]= 1599979481;
assign addr[45183]= 1649974225;
assign addr[45184]= 1697875851;
assign addr[45185]= 1743623590;
assign addr[45186]= 1787159411;
assign addr[45187]= 1828428082;
assign addr[45188]= 1867377253;
assign addr[45189]= 1903957513;
assign addr[45190]= 1938122457;
assign addr[45191]= 1969828744;
assign addr[45192]= 1999036154;
assign addr[45193]= 2025707632;
assign addr[45194]= 2049809346;
assign addr[45195]= 2071310720;
assign addr[45196]= 2090184478;
assign addr[45197]= 2106406677;
assign addr[45198]= 2119956737;
assign addr[45199]= 2130817471;
assign addr[45200]= 2138975100;
assign addr[45201]= 2144419275;
assign addr[45202]= 2147143090;
assign addr[45203]= 2147143090;
assign addr[45204]= 2144419275;
assign addr[45205]= 2138975100;
assign addr[45206]= 2130817471;
assign addr[45207]= 2119956737;
assign addr[45208]= 2106406677;
assign addr[45209]= 2090184478;
assign addr[45210]= 2071310720;
assign addr[45211]= 2049809346;
assign addr[45212]= 2025707632;
assign addr[45213]= 1999036154;
assign addr[45214]= 1969828744;
assign addr[45215]= 1938122457;
assign addr[45216]= 1903957513;
assign addr[45217]= 1867377253;
assign addr[45218]= 1828428082;
assign addr[45219]= 1787159411;
assign addr[45220]= 1743623590;
assign addr[45221]= 1697875851;
assign addr[45222]= 1649974225;
assign addr[45223]= 1599979481;
assign addr[45224]= 1547955041;
assign addr[45225]= 1493966902;
assign addr[45226]= 1438083551;
assign addr[45227]= 1380375881;
assign addr[45228]= 1320917099;
assign addr[45229]= 1259782632;
assign addr[45230]= 1197050035;
assign addr[45231]= 1132798888;
assign addr[45232]= 1067110699;
assign addr[45233]= 1000068799;
assign addr[45234]= 931758235;
assign addr[45235]= 862265664;
assign addr[45236]= 791679244;
assign addr[45237]= 720088517;
assign addr[45238]= 647584304;
assign addr[45239]= 574258580;
assign addr[45240]= 500204365;
assign addr[45241]= 425515602;
assign addr[45242]= 350287041;
assign addr[45243]= 274614114;
assign addr[45244]= 198592817;
assign addr[45245]= 122319591;
assign addr[45246]= 45891193;
assign addr[45247]= -30595422;
assign addr[45248]= -107043224;
assign addr[45249]= -183355234;
assign addr[45250]= -259434643;
assign addr[45251]= -335184940;
assign addr[45252]= -410510029;
assign addr[45253]= -485314355;
assign addr[45254]= -559503022;
assign addr[45255]= -632981917;
assign addr[45256]= -705657826;
assign addr[45257]= -777438554;
assign addr[45258]= -848233042;
assign addr[45259]= -917951481;
assign addr[45260]= -986505429;
assign addr[45261]= -1053807919;
assign addr[45262]= -1119773573;
assign addr[45263]= -1184318708;
assign addr[45264]= -1247361445;
assign addr[45265]= -1308821808;
assign addr[45266]= -1368621831;
assign addr[45267]= -1426685652;
assign addr[45268]= -1482939614;
assign addr[45269]= -1537312353;
assign addr[45270]= -1589734894;
assign addr[45271]= -1640140734;
assign addr[45272]= -1688465931;
assign addr[45273]= -1734649179;
assign addr[45274]= -1778631892;
assign addr[45275]= -1820358275;
assign addr[45276]= -1859775393;
assign addr[45277]= -1896833245;
assign addr[45278]= -1931484818;
assign addr[45279]= -1963686155;
assign addr[45280]= -1993396407;
assign addr[45281]= -2020577882;
assign addr[45282]= -2045196100;
assign addr[45283]= -2067219829;
assign addr[45284]= -2086621133;
assign addr[45285]= -2103375398;
assign addr[45286]= -2117461370;
assign addr[45287]= -2128861181;
assign addr[45288]= -2137560369;
assign addr[45289]= -2143547897;
assign addr[45290]= -2146816171;
assign addr[45291]= -2147361045;
assign addr[45292]= -2145181827;
assign addr[45293]= -2140281282;
assign addr[45294]= -2132665626;
assign addr[45295]= -2122344521;
assign addr[45296]= -2109331059;
assign addr[45297]= -2093641749;
assign addr[45298]= -2075296495;
assign addr[45299]= -2054318569;
assign addr[45300]= -2030734582;
assign addr[45301]= -2004574453;
assign addr[45302]= -1975871368;
assign addr[45303]= -1944661739;
assign addr[45304]= -1910985158;
assign addr[45305]= -1874884346;
assign addr[45306]= -1836405100;
assign addr[45307]= -1795596234;
assign addr[45308]= -1752509516;
assign addr[45309]= -1707199606;
assign addr[45310]= -1659723983;
assign addr[45311]= -1610142873;
assign addr[45312]= -1558519173;
assign addr[45313]= -1504918373;
assign addr[45314]= -1449408469;
assign addr[45315]= -1392059879;
assign addr[45316]= -1332945355;
assign addr[45317]= -1272139887;
assign addr[45318]= -1209720613;
assign addr[45319]= -1145766716;
assign addr[45320]= -1080359326;
assign addr[45321]= -1013581418;
assign addr[45322]= -945517704;
assign addr[45323]= -876254528;
assign addr[45324]= -805879757;
assign addr[45325]= -734482665;
assign addr[45326]= -662153826;
assign addr[45327]= -588984994;
assign addr[45328]= -515068990;
assign addr[45329]= -440499581;
assign addr[45330]= -365371365;
assign addr[45331]= -289779648;
assign addr[45332]= -213820322;
assign addr[45333]= -137589750;
assign addr[45334]= -61184634;
assign addr[45335]= 15298099;
assign addr[45336]= 91761426;
assign addr[45337]= 168108346;
assign addr[45338]= 244242007;
assign addr[45339]= 320065829;
assign addr[45340]= 395483624;
assign addr[45341]= 470399716;
assign addr[45342]= 544719071;
assign addr[45343]= 618347408;
assign addr[45344]= 691191324;
assign addr[45345]= 763158411;
assign addr[45346]= 834157373;
assign addr[45347]= 904098143;
assign addr[45348]= 972891995;
assign addr[45349]= 1040451659;
assign addr[45350]= 1106691431;
assign addr[45351]= 1171527280;
assign addr[45352]= 1234876957;
assign addr[45353]= 1296660098;
assign addr[45354]= 1356798326;
assign addr[45355]= 1415215352;
assign addr[45356]= 1471837070;
assign addr[45357]= 1526591649;
assign addr[45358]= 1579409630;
assign addr[45359]= 1630224009;
assign addr[45360]= 1678970324;
assign addr[45361]= 1725586737;
assign addr[45362]= 1770014111;
assign addr[45363]= 1812196087;
assign addr[45364]= 1852079154;
assign addr[45365]= 1889612716;
assign addr[45366]= 1924749160;
assign addr[45367]= 1957443913;
assign addr[45368]= 1987655498;
assign addr[45369]= 2015345591;
assign addr[45370]= 2040479063;
assign addr[45371]= 2063024031;
assign addr[45372]= 2082951896;
assign addr[45373]= 2100237377;
assign addr[45374]= 2114858546;
assign addr[45375]= 2126796855;
assign addr[45376]= 2136037160;
assign addr[45377]= 2142567738;
assign addr[45378]= 2146380306;
assign addr[45379]= 2147470025;
assign addr[45380]= 2145835515;
assign addr[45381]= 2141478848;
assign addr[45382]= 2134405552;
assign addr[45383]= 2124624598;
assign addr[45384]= 2112148396;
assign addr[45385]= 2096992772;
assign addr[45386]= 2079176953;
assign addr[45387]= 2058723538;
assign addr[45388]= 2035658475;
assign addr[45389]= 2010011024;
assign addr[45390]= 1981813720;
assign addr[45391]= 1951102334;
assign addr[45392]= 1917915825;
assign addr[45393]= 1882296293;
assign addr[45394]= 1844288924;
assign addr[45395]= 1803941934;
assign addr[45396]= 1761306505;
assign addr[45397]= 1716436725;
assign addr[45398]= 1669389513;
assign addr[45399]= 1620224553;
assign addr[45400]= 1569004214;
assign addr[45401]= 1515793473;
assign addr[45402]= 1460659832;
assign addr[45403]= 1403673233;
assign addr[45404]= 1344905966;
assign addr[45405]= 1284432584;
assign addr[45406]= 1222329801;
assign addr[45407]= 1158676398;
assign addr[45408]= 1093553126;
assign addr[45409]= 1027042599;
assign addr[45410]= 959229189;
assign addr[45411]= 890198924;
assign addr[45412]= 820039373;
assign addr[45413]= 748839539;
assign addr[45414]= 676689746;
assign addr[45415]= 603681519;
assign addr[45416]= 529907477;
assign addr[45417]= 455461206;
assign addr[45418]= 380437148;
assign addr[45419]= 304930476;
assign addr[45420]= 229036977;
assign addr[45421]= 152852926;
assign addr[45422]= 76474970;
assign addr[45423]= 0;
assign addr[45424]= -76474970;
assign addr[45425]= -152852926;
assign addr[45426]= -229036977;
assign addr[45427]= -304930476;
assign addr[45428]= -380437148;
assign addr[45429]= -455461206;
assign addr[45430]= -529907477;
assign addr[45431]= -603681519;
assign addr[45432]= -676689746;
assign addr[45433]= -748839539;
assign addr[45434]= -820039373;
assign addr[45435]= -890198924;
assign addr[45436]= -959229189;
assign addr[45437]= -1027042599;
assign addr[45438]= -1093553126;
assign addr[45439]= -1158676398;
assign addr[45440]= -1222329801;
assign addr[45441]= -1284432584;
assign addr[45442]= -1344905966;
assign addr[45443]= -1403673233;
assign addr[45444]= -1460659832;
assign addr[45445]= -1515793473;
assign addr[45446]= -1569004214;
assign addr[45447]= -1620224553;
assign addr[45448]= -1669389513;
assign addr[45449]= -1716436725;
assign addr[45450]= -1761306505;
assign addr[45451]= -1803941934;
assign addr[45452]= -1844288924;
assign addr[45453]= -1882296293;
assign addr[45454]= -1917915825;
assign addr[45455]= -1951102334;
assign addr[45456]= -1981813720;
assign addr[45457]= -2010011024;
assign addr[45458]= -2035658475;
assign addr[45459]= -2058723538;
assign addr[45460]= -2079176953;
assign addr[45461]= -2096992772;
assign addr[45462]= -2112148396;
assign addr[45463]= -2124624598;
assign addr[45464]= -2134405552;
assign addr[45465]= -2141478848;
assign addr[45466]= -2145835515;
assign addr[45467]= -2147470025;
assign addr[45468]= -2146380306;
assign addr[45469]= -2142567738;
assign addr[45470]= -2136037160;
assign addr[45471]= -2126796855;
assign addr[45472]= -2114858546;
assign addr[45473]= -2100237377;
assign addr[45474]= -2082951896;
assign addr[45475]= -2063024031;
assign addr[45476]= -2040479063;
assign addr[45477]= -2015345591;
assign addr[45478]= -1987655498;
assign addr[45479]= -1957443913;
assign addr[45480]= -1924749160;
assign addr[45481]= -1889612716;
assign addr[45482]= -1852079154;
assign addr[45483]= -1812196087;
assign addr[45484]= -1770014111;
assign addr[45485]= -1725586737;
assign addr[45486]= -1678970324;
assign addr[45487]= -1630224009;
assign addr[45488]= -1579409630;
assign addr[45489]= -1526591649;
assign addr[45490]= -1471837070;
assign addr[45491]= -1415215352;
assign addr[45492]= -1356798326;
assign addr[45493]= -1296660098;
assign addr[45494]= -1234876957;
assign addr[45495]= -1171527280;
assign addr[45496]= -1106691431;
assign addr[45497]= -1040451659;
assign addr[45498]= -972891995;
assign addr[45499]= -904098143;
assign addr[45500]= -834157373;
assign addr[45501]= -763158411;
assign addr[45502]= -691191324;
assign addr[45503]= -618347408;
assign addr[45504]= -544719071;
assign addr[45505]= -470399716;
assign addr[45506]= -395483624;
assign addr[45507]= -320065829;
assign addr[45508]= -244242007;
assign addr[45509]= -168108346;
assign addr[45510]= -91761426;
assign addr[45511]= -15298099;
assign addr[45512]= 61184634;
assign addr[45513]= 137589750;
assign addr[45514]= 213820322;
assign addr[45515]= 289779648;
assign addr[45516]= 365371365;
assign addr[45517]= 440499581;
assign addr[45518]= 515068990;
assign addr[45519]= 588984994;
assign addr[45520]= 662153826;
assign addr[45521]= 734482665;
assign addr[45522]= 805879757;
assign addr[45523]= 876254528;
assign addr[45524]= 945517704;
assign addr[45525]= 1013581418;
assign addr[45526]= 1080359326;
assign addr[45527]= 1145766716;
assign addr[45528]= 1209720613;
assign addr[45529]= 1272139887;
assign addr[45530]= 1332945355;
assign addr[45531]= 1392059879;
assign addr[45532]= 1449408469;
assign addr[45533]= 1504918373;
assign addr[45534]= 1558519173;
assign addr[45535]= 1610142873;
assign addr[45536]= 1659723983;
assign addr[45537]= 1707199606;
assign addr[45538]= 1752509516;
assign addr[45539]= 1795596234;
assign addr[45540]= 1836405100;
assign addr[45541]= 1874884346;
assign addr[45542]= 1910985158;
assign addr[45543]= 1944661739;
assign addr[45544]= 1975871368;
assign addr[45545]= 2004574453;
assign addr[45546]= 2030734582;
assign addr[45547]= 2054318569;
assign addr[45548]= 2075296495;
assign addr[45549]= 2093641749;
assign addr[45550]= 2109331059;
assign addr[45551]= 2122344521;
assign addr[45552]= 2132665626;
assign addr[45553]= 2140281282;
assign addr[45554]= 2145181827;
assign addr[45555]= 2147361045;
assign addr[45556]= 2146816171;
assign addr[45557]= 2143547897;
assign addr[45558]= 2137560369;
assign addr[45559]= 2128861181;
assign addr[45560]= 2117461370;
assign addr[45561]= 2103375398;
assign addr[45562]= 2086621133;
assign addr[45563]= 2067219829;
assign addr[45564]= 2045196100;
assign addr[45565]= 2020577882;
assign addr[45566]= 1993396407;
assign addr[45567]= 1963686155;
assign addr[45568]= 1931484818;
assign addr[45569]= 1896833245;
assign addr[45570]= 1859775393;
assign addr[45571]= 1820358275;
assign addr[45572]= 1778631892;
assign addr[45573]= 1734649179;
assign addr[45574]= 1688465931;
assign addr[45575]= 1640140734;
assign addr[45576]= 1589734894;
assign addr[45577]= 1537312353;
assign addr[45578]= 1482939614;
assign addr[45579]= 1426685652;
assign addr[45580]= 1368621831;
assign addr[45581]= 1308821808;
assign addr[45582]= 1247361445;
assign addr[45583]= 1184318708;
assign addr[45584]= 1119773573;
assign addr[45585]= 1053807919;
assign addr[45586]= 986505429;
assign addr[45587]= 917951481;
assign addr[45588]= 848233042;
assign addr[45589]= 777438554;
assign addr[45590]= 705657826;
assign addr[45591]= 632981917;
assign addr[45592]= 559503022;
assign addr[45593]= 485314355;
assign addr[45594]= 410510029;
assign addr[45595]= 335184940;
assign addr[45596]= 259434643;
assign addr[45597]= 183355234;
assign addr[45598]= 107043224;
assign addr[45599]= 30595422;
assign addr[45600]= -45891193;
assign addr[45601]= -122319591;
assign addr[45602]= -198592817;
assign addr[45603]= -274614114;
assign addr[45604]= -350287041;
assign addr[45605]= -425515602;
assign addr[45606]= -500204365;
assign addr[45607]= -574258580;
assign addr[45608]= -647584304;
assign addr[45609]= -720088517;
assign addr[45610]= -791679244;
assign addr[45611]= -862265664;
assign addr[45612]= -931758235;
assign addr[45613]= -1000068799;
assign addr[45614]= -1067110699;
assign addr[45615]= -1132798888;
assign addr[45616]= -1197050035;
assign addr[45617]= -1259782632;
assign addr[45618]= -1320917099;
assign addr[45619]= -1380375881;
assign addr[45620]= -1438083551;
assign addr[45621]= -1493966902;
assign addr[45622]= -1547955041;
assign addr[45623]= -1599979481;
assign addr[45624]= -1649974225;
assign addr[45625]= -1697875851;
assign addr[45626]= -1743623590;
assign addr[45627]= -1787159411;
assign addr[45628]= -1828428082;
assign addr[45629]= -1867377253;
assign addr[45630]= -1903957513;
assign addr[45631]= -1938122457;
assign addr[45632]= -1969828744;
assign addr[45633]= -1999036154;
assign addr[45634]= -2025707632;
assign addr[45635]= -2049809346;
assign addr[45636]= -2071310720;
assign addr[45637]= -2090184478;
assign addr[45638]= -2106406677;
assign addr[45639]= -2119956737;
assign addr[45640]= -2130817471;
assign addr[45641]= -2138975100;
assign addr[45642]= -2144419275;
assign addr[45643]= -2147143090;
assign addr[45644]= -2147143090;
assign addr[45645]= -2144419275;
assign addr[45646]= -2138975100;
assign addr[45647]= -2130817471;
assign addr[45648]= -2119956737;
assign addr[45649]= -2106406677;
assign addr[45650]= -2090184478;
assign addr[45651]= -2071310720;
assign addr[45652]= -2049809346;
assign addr[45653]= -2025707632;
assign addr[45654]= -1999036154;
assign addr[45655]= -1969828744;
assign addr[45656]= -1938122457;
assign addr[45657]= -1903957513;
assign addr[45658]= -1867377253;
assign addr[45659]= -1828428082;
assign addr[45660]= -1787159411;
assign addr[45661]= -1743623590;
assign addr[45662]= -1697875851;
assign addr[45663]= -1649974225;
assign addr[45664]= -1599979481;
assign addr[45665]= -1547955041;
assign addr[45666]= -1493966902;
assign addr[45667]= -1438083551;
assign addr[45668]= -1380375881;
assign addr[45669]= -1320917099;
assign addr[45670]= -1259782632;
assign addr[45671]= -1197050035;
assign addr[45672]= -1132798888;
assign addr[45673]= -1067110699;
assign addr[45674]= -1000068799;
assign addr[45675]= -931758235;
assign addr[45676]= -862265664;
assign addr[45677]= -791679244;
assign addr[45678]= -720088517;
assign addr[45679]= -647584304;
assign addr[45680]= -574258580;
assign addr[45681]= -500204365;
assign addr[45682]= -425515602;
assign addr[45683]= -350287041;
assign addr[45684]= -274614114;
assign addr[45685]= -198592817;
assign addr[45686]= -122319591;
assign addr[45687]= -45891193;
assign addr[45688]= 30595422;
assign addr[45689]= 107043224;
assign addr[45690]= 183355234;
assign addr[45691]= 259434643;
assign addr[45692]= 335184940;
assign addr[45693]= 410510029;
assign addr[45694]= 485314355;
assign addr[45695]= 559503022;
assign addr[45696]= 632981917;
assign addr[45697]= 705657826;
assign addr[45698]= 777438554;
assign addr[45699]= 848233042;
assign addr[45700]= 917951481;
assign addr[45701]= 986505429;
assign addr[45702]= 1053807919;
assign addr[45703]= 1119773573;
assign addr[45704]= 1184318708;
assign addr[45705]= 1247361445;
assign addr[45706]= 1308821808;
assign addr[45707]= 1368621831;
assign addr[45708]= 1426685652;
assign addr[45709]= 1482939614;
assign addr[45710]= 1537312353;
assign addr[45711]= 1589734894;
assign addr[45712]= 1640140734;
assign addr[45713]= 1688465931;
assign addr[45714]= 1734649179;
assign addr[45715]= 1778631892;
assign addr[45716]= 1820358275;
assign addr[45717]= 1859775393;
assign addr[45718]= 1896833245;
assign addr[45719]= 1931484818;
assign addr[45720]= 1963686155;
assign addr[45721]= 1993396407;
assign addr[45722]= 2020577882;
assign addr[45723]= 2045196100;
assign addr[45724]= 2067219829;
assign addr[45725]= 2086621133;
assign addr[45726]= 2103375398;
assign addr[45727]= 2117461370;
assign addr[45728]= 2128861181;
assign addr[45729]= 2137560369;
assign addr[45730]= 2143547897;
assign addr[45731]= 2146816171;
assign addr[45732]= 2147361045;
assign addr[45733]= 2145181827;
assign addr[45734]= 2140281282;
assign addr[45735]= 2132665626;
assign addr[45736]= 2122344521;
assign addr[45737]= 2109331059;
assign addr[45738]= 2093641749;
assign addr[45739]= 2075296495;
assign addr[45740]= 2054318569;
assign addr[45741]= 2030734582;
assign addr[45742]= 2004574453;
assign addr[45743]= 1975871368;
assign addr[45744]= 1944661739;
assign addr[45745]= 1910985158;
assign addr[45746]= 1874884346;
assign addr[45747]= 1836405100;
assign addr[45748]= 1795596234;
assign addr[45749]= 1752509516;
assign addr[45750]= 1707199606;
assign addr[45751]= 1659723983;
assign addr[45752]= 1610142873;
assign addr[45753]= 1558519173;
assign addr[45754]= 1504918373;
assign addr[45755]= 1449408469;
assign addr[45756]= 1392059879;
assign addr[45757]= 1332945355;
assign addr[45758]= 1272139887;
assign addr[45759]= 1209720613;
assign addr[45760]= 1145766716;
assign addr[45761]= 1080359326;
assign addr[45762]= 1013581418;
assign addr[45763]= 945517704;
assign addr[45764]= 876254528;
assign addr[45765]= 805879757;
assign addr[45766]= 734482665;
assign addr[45767]= 662153826;
assign addr[45768]= 588984994;
assign addr[45769]= 515068990;
assign addr[45770]= 440499581;
assign addr[45771]= 365371365;
assign addr[45772]= 289779648;
assign addr[45773]= 213820322;
assign addr[45774]= 137589750;
assign addr[45775]= 61184634;
assign addr[45776]= -15298099;
assign addr[45777]= -91761426;
assign addr[45778]= -168108346;
assign addr[45779]= -244242007;
assign addr[45780]= -320065829;
assign addr[45781]= -395483624;
assign addr[45782]= -470399716;
assign addr[45783]= -544719071;
assign addr[45784]= -618347408;
assign addr[45785]= -691191324;
assign addr[45786]= -763158411;
assign addr[45787]= -834157373;
assign addr[45788]= -904098143;
assign addr[45789]= -972891995;
assign addr[45790]= -1040451659;
assign addr[45791]= -1106691431;
assign addr[45792]= -1171527280;
assign addr[45793]= -1234876957;
assign addr[45794]= -1296660098;
assign addr[45795]= -1356798326;
assign addr[45796]= -1415215352;
assign addr[45797]= -1471837070;
assign addr[45798]= -1526591649;
assign addr[45799]= -1579409630;
assign addr[45800]= -1630224009;
assign addr[45801]= -1678970324;
assign addr[45802]= -1725586737;
assign addr[45803]= -1770014111;
assign addr[45804]= -1812196087;
assign addr[45805]= -1852079154;
assign addr[45806]= -1889612716;
assign addr[45807]= -1924749160;
assign addr[45808]= -1957443913;
assign addr[45809]= -1987655498;
assign addr[45810]= -2015345591;
assign addr[45811]= -2040479063;
assign addr[45812]= -2063024031;
assign addr[45813]= -2082951896;
assign addr[45814]= -2100237377;
assign addr[45815]= -2114858546;
assign addr[45816]= -2126796855;
assign addr[45817]= -2136037160;
assign addr[45818]= -2142567738;
assign addr[45819]= -2146380306;
assign addr[45820]= -2147470025;
assign addr[45821]= -2145835515;
assign addr[45822]= -2141478848;
assign addr[45823]= -2134405552;
assign addr[45824]= -2124624598;
assign addr[45825]= -2112148396;
assign addr[45826]= -2096992772;
assign addr[45827]= -2079176953;
assign addr[45828]= -2058723538;
assign addr[45829]= -2035658475;
assign addr[45830]= -2010011024;
assign addr[45831]= -1981813720;
assign addr[45832]= -1951102334;
assign addr[45833]= -1917915825;
assign addr[45834]= -1882296293;
assign addr[45835]= -1844288924;
assign addr[45836]= -1803941934;
assign addr[45837]= -1761306505;
assign addr[45838]= -1716436725;
assign addr[45839]= -1669389513;
assign addr[45840]= -1620224553;
assign addr[45841]= -1569004214;
assign addr[45842]= -1515793473;
assign addr[45843]= -1460659832;
assign addr[45844]= -1403673233;
assign addr[45845]= -1344905966;
assign addr[45846]= -1284432584;
assign addr[45847]= -1222329801;
assign addr[45848]= -1158676398;
assign addr[45849]= -1093553126;
assign addr[45850]= -1027042599;
assign addr[45851]= -959229189;
assign addr[45852]= -890198924;
assign addr[45853]= -820039373;
assign addr[45854]= -748839539;
assign addr[45855]= -676689746;
assign addr[45856]= -603681519;
assign addr[45857]= -529907477;
assign addr[45858]= -455461206;
assign addr[45859]= -380437148;
assign addr[45860]= -304930476;
assign addr[45861]= -229036977;
assign addr[45862]= -152852926;
assign addr[45863]= -76474970;
assign addr[45864]= 0;
assign addr[45865]= 76474970;
assign addr[45866]= 152852926;
assign addr[45867]= 229036977;
assign addr[45868]= 304930476;
assign addr[45869]= 380437148;
assign addr[45870]= 455461206;
assign addr[45871]= 529907477;
assign addr[45872]= 603681519;
assign addr[45873]= 676689746;
assign addr[45874]= 748839539;
assign addr[45875]= 820039373;
assign addr[45876]= 890198924;
assign addr[45877]= 959229189;
assign addr[45878]= 1027042599;
assign addr[45879]= 1093553126;
assign addr[45880]= 1158676398;
assign addr[45881]= 1222329801;
assign addr[45882]= 1284432584;
assign addr[45883]= 1344905966;
assign addr[45884]= 1403673233;
assign addr[45885]= 1460659832;
assign addr[45886]= 1515793473;
assign addr[45887]= 1569004214;
assign addr[45888]= 1620224553;
assign addr[45889]= 1669389513;
assign addr[45890]= 1716436725;
assign addr[45891]= 1761306505;
assign addr[45892]= 1803941934;
assign addr[45893]= 1844288924;
assign addr[45894]= 1882296293;
assign addr[45895]= 1917915825;
assign addr[45896]= 1951102334;
assign addr[45897]= 1981813720;
assign addr[45898]= 2010011024;
assign addr[45899]= 2035658475;
assign addr[45900]= 2058723538;
assign addr[45901]= 2079176953;
assign addr[45902]= 2096992772;
assign addr[45903]= 2112148396;
assign addr[45904]= 2124624598;
assign addr[45905]= 2134405552;
assign addr[45906]= 2141478848;
assign addr[45907]= 2145835515;
assign addr[45908]= 2147470025;
assign addr[45909]= 2146380306;
assign addr[45910]= 2142567738;
assign addr[45911]= 2136037160;
assign addr[45912]= 2126796855;
assign addr[45913]= 2114858546;
assign addr[45914]= 2100237377;
assign addr[45915]= 2082951896;
assign addr[45916]= 2063024031;
assign addr[45917]= 2040479063;
assign addr[45918]= 2015345591;
assign addr[45919]= 1987655498;
assign addr[45920]= 1957443913;
assign addr[45921]= 1924749160;
assign addr[45922]= 1889612716;
assign addr[45923]= 1852079154;
assign addr[45924]= 1812196087;
assign addr[45925]= 1770014111;
assign addr[45926]= 1725586737;
assign addr[45927]= 1678970324;
assign addr[45928]= 1630224009;
assign addr[45929]= 1579409630;
assign addr[45930]= 1526591649;
assign addr[45931]= 1471837070;
assign addr[45932]= 1415215352;
assign addr[45933]= 1356798326;
assign addr[45934]= 1296660098;
assign addr[45935]= 1234876957;
assign addr[45936]= 1171527280;
assign addr[45937]= 1106691431;
assign addr[45938]= 1040451659;
assign addr[45939]= 972891995;
assign addr[45940]= 904098143;
assign addr[45941]= 834157373;
assign addr[45942]= 763158411;
assign addr[45943]= 691191324;
assign addr[45944]= 618347408;
assign addr[45945]= 544719071;
assign addr[45946]= 470399716;
assign addr[45947]= 395483624;
assign addr[45948]= 320065829;
assign addr[45949]= 244242007;
assign addr[45950]= 168108346;
assign addr[45951]= 91761426;
assign addr[45952]= 15298099;
assign addr[45953]= -61184634;
assign addr[45954]= -137589750;
assign addr[45955]= -213820322;
assign addr[45956]= -289779648;
assign addr[45957]= -365371365;
assign addr[45958]= -440499581;
assign addr[45959]= -515068990;
assign addr[45960]= -588984994;
assign addr[45961]= -662153826;
assign addr[45962]= -734482665;
assign addr[45963]= -805879757;
assign addr[45964]= -876254528;
assign addr[45965]= -945517704;
assign addr[45966]= -1013581418;
assign addr[45967]= -1080359326;
assign addr[45968]= -1145766716;
assign addr[45969]= -1209720613;
assign addr[45970]= -1272139887;
assign addr[45971]= -1332945355;
assign addr[45972]= -1392059879;
assign addr[45973]= -1449408469;
assign addr[45974]= -1504918373;
assign addr[45975]= -1558519173;
assign addr[45976]= -1610142873;
assign addr[45977]= -1659723983;
assign addr[45978]= -1707199606;
assign addr[45979]= -1752509516;
assign addr[45980]= -1795596234;
assign addr[45981]= -1836405100;
assign addr[45982]= -1874884346;
assign addr[45983]= -1910985158;
assign addr[45984]= -1944661739;
assign addr[45985]= -1975871368;
assign addr[45986]= -2004574453;
assign addr[45987]= -2030734582;
assign addr[45988]= -2054318569;
assign addr[45989]= -2075296495;
assign addr[45990]= -2093641749;
assign addr[45991]= -2109331059;
assign addr[45992]= -2122344521;
assign addr[45993]= -2132665626;
assign addr[45994]= -2140281282;
assign addr[45995]= -2145181827;
assign addr[45996]= -2147361045;
assign addr[45997]= -2146816171;
assign addr[45998]= -2143547897;
assign addr[45999]= -2137560369;
assign addr[46000]= -2128861181;
assign addr[46001]= -2117461370;
assign addr[46002]= -2103375398;
assign addr[46003]= -2086621133;
assign addr[46004]= -2067219829;
assign addr[46005]= -2045196100;
assign addr[46006]= -2020577882;
assign addr[46007]= -1993396407;
assign addr[46008]= -1963686155;
assign addr[46009]= -1931484818;
assign addr[46010]= -1896833245;
assign addr[46011]= -1859775393;
assign addr[46012]= -1820358275;
assign addr[46013]= -1778631892;
assign addr[46014]= -1734649179;
assign addr[46015]= -1688465931;
assign addr[46016]= -1640140734;
assign addr[46017]= -1589734894;
assign addr[46018]= -1537312353;
assign addr[46019]= -1482939614;
assign addr[46020]= -1426685652;
assign addr[46021]= -1368621831;
assign addr[46022]= -1308821808;
assign addr[46023]= -1247361445;
assign addr[46024]= -1184318708;
assign addr[46025]= -1119773573;
assign addr[46026]= -1053807919;
assign addr[46027]= -986505429;
assign addr[46028]= -917951481;
assign addr[46029]= -848233042;
assign addr[46030]= -777438554;
assign addr[46031]= -705657826;
assign addr[46032]= -632981917;
assign addr[46033]= -559503022;
assign addr[46034]= -485314355;
assign addr[46035]= -410510029;
assign addr[46036]= -335184940;
assign addr[46037]= -259434643;
assign addr[46038]= -183355234;
assign addr[46039]= -107043224;
assign addr[46040]= -30595422;
assign addr[46041]= 45891193;
assign addr[46042]= 122319591;
assign addr[46043]= 198592817;
assign addr[46044]= 274614114;
assign addr[46045]= 350287041;
assign addr[46046]= 425515602;
assign addr[46047]= 500204365;
assign addr[46048]= 574258580;
assign addr[46049]= 647584304;
assign addr[46050]= 720088517;
assign addr[46051]= 791679244;
assign addr[46052]= 862265664;
assign addr[46053]= 931758235;
assign addr[46054]= 1000068799;
assign addr[46055]= 1067110699;
assign addr[46056]= 1132798888;
assign addr[46057]= 1197050035;
assign addr[46058]= 1259782632;
assign addr[46059]= 1320917099;
assign addr[46060]= 1380375881;
assign addr[46061]= 1438083551;
assign addr[46062]= 1493966902;
assign addr[46063]= 1547955041;
assign addr[46064]= 1599979481;
assign addr[46065]= 1649974225;
assign addr[46066]= 1697875851;
assign addr[46067]= 1743623590;
assign addr[46068]= 1787159411;
assign addr[46069]= 1828428082;
assign addr[46070]= 1867377253;
assign addr[46071]= 1903957513;
assign addr[46072]= 1938122457;
assign addr[46073]= 1969828744;
assign addr[46074]= 1999036154;
assign addr[46075]= 2025707632;
assign addr[46076]= 2049809346;
assign addr[46077]= 2071310720;
assign addr[46078]= 2090184478;
assign addr[46079]= 2106406677;
assign addr[46080]= 2119956737;
assign addr[46081]= 2130817471;
assign addr[46082]= 2138975100;
assign addr[46083]= 2144419275;
assign addr[46084]= 2147143090;
assign addr[46085]= 2147143090;
assign addr[46086]= 2144419275;
assign addr[46087]= 2138975100;
assign addr[46088]= 2130817471;
assign addr[46089]= 2119956737;
assign addr[46090]= 2106406677;
assign addr[46091]= 2090184478;
assign addr[46092]= 2071310720;
assign addr[46093]= 2049809346;
assign addr[46094]= 2025707632;
assign addr[46095]= 1999036154;
assign addr[46096]= 1969828744;
assign addr[46097]= 1938122457;
assign addr[46098]= 1903957513;
assign addr[46099]= 1867377253;
assign addr[46100]= 1828428082;
assign addr[46101]= 1787159411;
assign addr[46102]= 1743623590;
assign addr[46103]= 1697875851;
assign addr[46104]= 1649974225;
assign addr[46105]= 1599979481;
assign addr[46106]= 1547955041;
assign addr[46107]= 1493966902;
assign addr[46108]= 1438083551;
assign addr[46109]= 1380375881;
assign addr[46110]= 1320917099;
assign addr[46111]= 1259782632;
assign addr[46112]= 1197050035;
assign addr[46113]= 1132798888;
assign addr[46114]= 1067110699;
assign addr[46115]= 1000068799;
assign addr[46116]= 931758235;
assign addr[46117]= 862265664;
assign addr[46118]= 791679244;
assign addr[46119]= 720088517;
assign addr[46120]= 647584304;
assign addr[46121]= 574258580;
assign addr[46122]= 500204365;
assign addr[46123]= 425515602;
assign addr[46124]= 350287041;
assign addr[46125]= 274614114;
assign addr[46126]= 198592817;
assign addr[46127]= 122319591;
assign addr[46128]= 45891193;
assign addr[46129]= -30595422;
assign addr[46130]= -107043224;
assign addr[46131]= -183355234;
assign addr[46132]= -259434643;
assign addr[46133]= -335184940;
assign addr[46134]= -410510029;
assign addr[46135]= -485314355;
assign addr[46136]= -559503022;
assign addr[46137]= -632981917;
assign addr[46138]= -705657826;
assign addr[46139]= -777438554;
assign addr[46140]= -848233042;
assign addr[46141]= -917951481;
assign addr[46142]= -986505429;
assign addr[46143]= -1053807919;
assign addr[46144]= -1119773573;
assign addr[46145]= -1184318708;
assign addr[46146]= -1247361445;
assign addr[46147]= -1308821808;
assign addr[46148]= -1368621831;
assign addr[46149]= -1426685652;
assign addr[46150]= -1482939614;
assign addr[46151]= -1537312353;
assign addr[46152]= -1589734894;
assign addr[46153]= -1640140734;
assign addr[46154]= -1688465931;
assign addr[46155]= -1734649179;
assign addr[46156]= -1778631892;
assign addr[46157]= -1820358275;
assign addr[46158]= -1859775393;
assign addr[46159]= -1896833245;
assign addr[46160]= -1931484818;
assign addr[46161]= -1963686155;
assign addr[46162]= -1993396407;
assign addr[46163]= -2020577882;
assign addr[46164]= -2045196100;
assign addr[46165]= -2067219829;
assign addr[46166]= -2086621133;
assign addr[46167]= -2103375398;
assign addr[46168]= -2117461370;
assign addr[46169]= -2128861181;
assign addr[46170]= -2137560369;
assign addr[46171]= -2143547897;
assign addr[46172]= -2146816171;
assign addr[46173]= -2147361045;
assign addr[46174]= -2145181827;
assign addr[46175]= -2140281282;
assign addr[46176]= -2132665626;
assign addr[46177]= -2122344521;
assign addr[46178]= -2109331059;
assign addr[46179]= -2093641749;
assign addr[46180]= -2075296495;
assign addr[46181]= -2054318569;
assign addr[46182]= -2030734582;
assign addr[46183]= -2004574453;
assign addr[46184]= -1975871368;
assign addr[46185]= -1944661739;
assign addr[46186]= -1910985158;
assign addr[46187]= -1874884346;
assign addr[46188]= -1836405100;
assign addr[46189]= -1795596234;
assign addr[46190]= -1752509516;
assign addr[46191]= -1707199606;
assign addr[46192]= -1659723983;
assign addr[46193]= -1610142873;
assign addr[46194]= -1558519173;
assign addr[46195]= -1504918373;
assign addr[46196]= -1449408469;
assign addr[46197]= -1392059879;
assign addr[46198]= -1332945355;
assign addr[46199]= -1272139887;
assign addr[46200]= -1209720613;
assign addr[46201]= -1145766716;
assign addr[46202]= -1080359326;
assign addr[46203]= -1013581418;
assign addr[46204]= -945517704;
assign addr[46205]= -876254528;
assign addr[46206]= -805879757;
assign addr[46207]= -734482665;
assign addr[46208]= -662153826;
assign addr[46209]= -588984994;
assign addr[46210]= -515068990;
assign addr[46211]= -440499581;
assign addr[46212]= -365371365;
assign addr[46213]= -289779648;
assign addr[46214]= -213820322;
assign addr[46215]= -137589750;
assign addr[46216]= -61184634;
assign addr[46217]= 15298099;
assign addr[46218]= 91761426;
assign addr[46219]= 168108346;
assign addr[46220]= 244242007;
assign addr[46221]= 320065829;
assign addr[46222]= 395483624;
assign addr[46223]= 470399716;
assign addr[46224]= 544719071;
assign addr[46225]= 618347408;
assign addr[46226]= 691191324;
assign addr[46227]= 763158411;
assign addr[46228]= 834157373;
assign addr[46229]= 904098143;
assign addr[46230]= 972891995;
assign addr[46231]= 1040451659;
assign addr[46232]= 1106691431;
assign addr[46233]= 1171527280;
assign addr[46234]= 1234876957;
assign addr[46235]= 1296660098;
assign addr[46236]= 1356798326;
assign addr[46237]= 1415215352;
assign addr[46238]= 1471837070;
assign addr[46239]= 1526591649;
assign addr[46240]= 1579409630;
assign addr[46241]= 1630224009;
assign addr[46242]= 1678970324;
assign addr[46243]= 1725586737;
assign addr[46244]= 1770014111;
assign addr[46245]= 1812196087;
assign addr[46246]= 1852079154;
assign addr[46247]= 1889612716;
assign addr[46248]= 1924749160;
assign addr[46249]= 1957443913;
assign addr[46250]= 1987655498;
assign addr[46251]= 2015345591;
assign addr[46252]= 2040479063;
assign addr[46253]= 2063024031;
assign addr[46254]= 2082951896;
assign addr[46255]= 2100237377;
assign addr[46256]= 2114858546;
assign addr[46257]= 2126796855;
assign addr[46258]= 2136037160;
assign addr[46259]= 2142567738;
assign addr[46260]= 2146380306;
assign addr[46261]= 2147470025;
assign addr[46262]= 2145835515;
assign addr[46263]= 2141478848;
assign addr[46264]= 2134405552;
assign addr[46265]= 2124624598;
assign addr[46266]= 2112148396;
assign addr[46267]= 2096992772;
assign addr[46268]= 2079176953;
assign addr[46269]= 2058723538;
assign addr[46270]= 2035658475;
assign addr[46271]= 2010011024;
assign addr[46272]= 1981813720;
assign addr[46273]= 1951102334;
assign addr[46274]= 1917915825;
assign addr[46275]= 1882296293;
assign addr[46276]= 1844288924;
assign addr[46277]= 1803941934;
assign addr[46278]= 1761306505;
assign addr[46279]= 1716436725;
assign addr[46280]= 1669389513;
assign addr[46281]= 1620224553;
assign addr[46282]= 1569004214;
assign addr[46283]= 1515793473;
assign addr[46284]= 1460659832;
assign addr[46285]= 1403673233;
assign addr[46286]= 1344905966;
assign addr[46287]= 1284432584;
assign addr[46288]= 1222329801;
assign addr[46289]= 1158676398;
assign addr[46290]= 1093553126;
assign addr[46291]= 1027042599;
assign addr[46292]= 959229189;
assign addr[46293]= 890198924;
assign addr[46294]= 820039373;
assign addr[46295]= 748839539;
assign addr[46296]= 676689746;
assign addr[46297]= 603681519;
assign addr[46298]= 529907477;
assign addr[46299]= 455461206;
assign addr[46300]= 380437148;
assign addr[46301]= 304930476;
assign addr[46302]= 229036977;
assign addr[46303]= 152852926;
assign addr[46304]= 76474970;
assign addr[46305]= 0;
assign addr[46306]= -76474970;
assign addr[46307]= -152852926;
assign addr[46308]= -229036977;
assign addr[46309]= -304930476;
assign addr[46310]= -380437148;
assign addr[46311]= -455461206;
assign addr[46312]= -529907477;
assign addr[46313]= -603681519;
assign addr[46314]= -676689746;
assign addr[46315]= -748839539;
assign addr[46316]= -820039373;
assign addr[46317]= -890198924;
assign addr[46318]= -959229189;
assign addr[46319]= -1027042599;
assign addr[46320]= -1093553126;
assign addr[46321]= -1158676398;
assign addr[46322]= -1222329801;
assign addr[46323]= -1284432584;
assign addr[46324]= -1344905966;
assign addr[46325]= -1403673233;
assign addr[46326]= -1460659832;
assign addr[46327]= -1515793473;
assign addr[46328]= -1569004214;
assign addr[46329]= -1620224553;
assign addr[46330]= -1669389513;
assign addr[46331]= -1716436725;
assign addr[46332]= -1761306505;
assign addr[46333]= -1803941934;
assign addr[46334]= -1844288924;
assign addr[46335]= -1882296293;
assign addr[46336]= -1917915825;
assign addr[46337]= -1951102334;
assign addr[46338]= -1981813720;
assign addr[46339]= -2010011024;
assign addr[46340]= -2035658475;
assign addr[46341]= -2058723538;
assign addr[46342]= -2079176953;
assign addr[46343]= -2096992772;
assign addr[46344]= -2112148396;
assign addr[46345]= -2124624598;
assign addr[46346]= -2134405552;
assign addr[46347]= -2141478848;
assign addr[46348]= -2145835515;
assign addr[46349]= -2147470025;
assign addr[46350]= -2146380306;
assign addr[46351]= -2142567738;
assign addr[46352]= -2136037160;
assign addr[46353]= -2126796855;
assign addr[46354]= -2114858546;
assign addr[46355]= -2100237377;
assign addr[46356]= -2082951896;
assign addr[46357]= -2063024031;
assign addr[46358]= -2040479063;
assign addr[46359]= -2015345591;
assign addr[46360]= -1987655498;
assign addr[46361]= -1957443913;
assign addr[46362]= -1924749160;
assign addr[46363]= -1889612716;
assign addr[46364]= -1852079154;
assign addr[46365]= -1812196087;
assign addr[46366]= -1770014111;
assign addr[46367]= -1725586737;
assign addr[46368]= -1678970324;
assign addr[46369]= -1630224009;
assign addr[46370]= -1579409630;
assign addr[46371]= -1526591649;
assign addr[46372]= -1471837070;
assign addr[46373]= -1415215352;
assign addr[46374]= -1356798326;
assign addr[46375]= -1296660098;
assign addr[46376]= -1234876957;
assign addr[46377]= -1171527280;
assign addr[46378]= -1106691431;
assign addr[46379]= -1040451659;
assign addr[46380]= -972891995;
assign addr[46381]= -904098143;
assign addr[46382]= -834157373;
assign addr[46383]= -763158411;
assign addr[46384]= -691191324;
assign addr[46385]= -618347408;
assign addr[46386]= -544719071;
assign addr[46387]= -470399716;
assign addr[46388]= -395483624;
assign addr[46389]= -320065829;
assign addr[46390]= -244242007;
assign addr[46391]= -168108346;
assign addr[46392]= -91761426;
assign addr[46393]= -15298099;
assign addr[46394]= 61184634;
assign addr[46395]= 137589750;
assign addr[46396]= 213820322;
assign addr[46397]= 289779648;
assign addr[46398]= 365371365;
assign addr[46399]= 440499581;
assign addr[46400]= 515068990;
assign addr[46401]= 588984994;
assign addr[46402]= 662153826;
assign addr[46403]= 734482665;
assign addr[46404]= 805879757;
assign addr[46405]= 876254528;
assign addr[46406]= 945517704;
assign addr[46407]= 1013581418;
assign addr[46408]= 1080359326;
assign addr[46409]= 1145766716;
assign addr[46410]= 1209720613;
assign addr[46411]= 1272139887;
assign addr[46412]= 1332945355;
assign addr[46413]= 1392059879;
assign addr[46414]= 1449408469;
assign addr[46415]= 1504918373;
assign addr[46416]= 1558519173;
assign addr[46417]= 1610142873;
assign addr[46418]= 1659723983;
assign addr[46419]= 1707199606;
assign addr[46420]= 1752509516;
assign addr[46421]= 1795596234;
assign addr[46422]= 1836405100;
assign addr[46423]= 1874884346;
assign addr[46424]= 1910985158;
assign addr[46425]= 1944661739;
assign addr[46426]= 1975871368;
assign addr[46427]= 2004574453;
assign addr[46428]= 2030734582;
assign addr[46429]= 2054318569;
assign addr[46430]= 2075296495;
assign addr[46431]= 2093641749;
assign addr[46432]= 2109331059;
assign addr[46433]= 2122344521;
assign addr[46434]= 2132665626;
assign addr[46435]= 2140281282;
assign addr[46436]= 2145181827;
assign addr[46437]= 2147361045;
assign addr[46438]= 2146816171;
assign addr[46439]= 2143547897;
assign addr[46440]= 2137560369;
assign addr[46441]= 2128861181;
assign addr[46442]= 2117461370;
assign addr[46443]= 2103375398;
assign addr[46444]= 2086621133;
assign addr[46445]= 2067219829;
assign addr[46446]= 2045196100;
assign addr[46447]= 2020577882;
assign addr[46448]= 1993396407;
assign addr[46449]= 1963686155;
assign addr[46450]= 1931484818;
assign addr[46451]= 1896833245;
assign addr[46452]= 1859775393;
assign addr[46453]= 1820358275;
assign addr[46454]= 1778631892;
assign addr[46455]= 1734649179;
assign addr[46456]= 1688465931;
assign addr[46457]= 1640140734;
assign addr[46458]= 1589734894;
assign addr[46459]= 1537312353;
assign addr[46460]= 1482939614;
assign addr[46461]= 1426685652;
assign addr[46462]= 1368621831;
assign addr[46463]= 1308821808;
assign addr[46464]= 1247361445;
assign addr[46465]= 1184318708;
assign addr[46466]= 1119773573;
assign addr[46467]= 1053807919;
assign addr[46468]= 986505429;
assign addr[46469]= 917951481;
assign addr[46470]= 848233042;
assign addr[46471]= 777438554;
assign addr[46472]= 705657826;
assign addr[46473]= 632981917;
assign addr[46474]= 559503022;
assign addr[46475]= 485314355;
assign addr[46476]= 410510029;
assign addr[46477]= 335184940;
assign addr[46478]= 259434643;
assign addr[46479]= 183355234;
assign addr[46480]= 107043224;
assign addr[46481]= 30595422;
assign addr[46482]= -45891193;
assign addr[46483]= -122319591;
assign addr[46484]= -198592817;
assign addr[46485]= -274614114;
assign addr[46486]= -350287041;
assign addr[46487]= -425515602;
assign addr[46488]= -500204365;
assign addr[46489]= -574258580;
assign addr[46490]= -647584304;
assign addr[46491]= -720088517;
assign addr[46492]= -791679244;
assign addr[46493]= -862265664;
assign addr[46494]= -931758235;
assign addr[46495]= -1000068799;
assign addr[46496]= -1067110699;
assign addr[46497]= -1132798888;
assign addr[46498]= -1197050035;
assign addr[46499]= -1259782632;
assign addr[46500]= -1320917099;
assign addr[46501]= -1380375881;
assign addr[46502]= -1438083551;
assign addr[46503]= -1493966902;
assign addr[46504]= -1547955041;
assign addr[46505]= -1599979481;
assign addr[46506]= -1649974225;
assign addr[46507]= -1697875851;
assign addr[46508]= -1743623590;
assign addr[46509]= -1787159411;
assign addr[46510]= -1828428082;
assign addr[46511]= -1867377253;
assign addr[46512]= -1903957513;
assign addr[46513]= -1938122457;
assign addr[46514]= -1969828744;
assign addr[46515]= -1999036154;
assign addr[46516]= -2025707632;
assign addr[46517]= -2049809346;
assign addr[46518]= -2071310720;
assign addr[46519]= -2090184478;
assign addr[46520]= -2106406677;
assign addr[46521]= -2119956737;
assign addr[46522]= -2130817471;
assign addr[46523]= -2138975100;
assign addr[46524]= -2144419275;
assign addr[46525]= -2147143090;
assign addr[46526]= -2147143090;
assign addr[46527]= -2144419275;
assign addr[46528]= -2138975100;
assign addr[46529]= -2130817471;
assign addr[46530]= -2119956737;
assign addr[46531]= -2106406677;
assign addr[46532]= -2090184478;
assign addr[46533]= -2071310720;
assign addr[46534]= -2049809346;
assign addr[46535]= -2025707632;
assign addr[46536]= -1999036154;
assign addr[46537]= -1969828744;
assign addr[46538]= -1938122457;
assign addr[46539]= -1903957513;
assign addr[46540]= -1867377253;
assign addr[46541]= -1828428082;
assign addr[46542]= -1787159411;
assign addr[46543]= -1743623590;
assign addr[46544]= -1697875851;
assign addr[46545]= -1649974225;
assign addr[46546]= -1599979481;
assign addr[46547]= -1547955041;
assign addr[46548]= -1493966902;
assign addr[46549]= -1438083551;
assign addr[46550]= -1380375881;
assign addr[46551]= -1320917099;
assign addr[46552]= -1259782632;
assign addr[46553]= -1197050035;
assign addr[46554]= -1132798888;
assign addr[46555]= -1067110699;
assign addr[46556]= -1000068799;
assign addr[46557]= -931758235;
assign addr[46558]= -862265664;
assign addr[46559]= -791679244;
assign addr[46560]= -720088517;
assign addr[46561]= -647584304;
assign addr[46562]= -574258580;
assign addr[46563]= -500204365;
assign addr[46564]= -425515602;
assign addr[46565]= -350287041;
assign addr[46566]= -274614114;
assign addr[46567]= -198592817;
assign addr[46568]= -122319591;
assign addr[46569]= -45891193;
assign addr[46570]= 30595422;
assign addr[46571]= 107043224;
assign addr[46572]= 183355234;
assign addr[46573]= 259434643;
assign addr[46574]= 335184940;
assign addr[46575]= 410510029;
assign addr[46576]= 485314355;
assign addr[46577]= 559503022;
assign addr[46578]= 632981917;
assign addr[46579]= 705657826;
assign addr[46580]= 777438554;
assign addr[46581]= 848233042;
assign addr[46582]= 917951481;
assign addr[46583]= 986505429;
assign addr[46584]= 1053807919;
assign addr[46585]= 1119773573;
assign addr[46586]= 1184318708;
assign addr[46587]= 1247361445;
assign addr[46588]= 1308821808;
assign addr[46589]= 1368621831;
assign addr[46590]= 1426685652;
assign addr[46591]= 1482939614;
assign addr[46592]= 1537312353;
assign addr[46593]= 1589734894;
assign addr[46594]= 1640140734;
assign addr[46595]= 1688465931;
assign addr[46596]= 1734649179;
assign addr[46597]= 1778631892;
assign addr[46598]= 1820358275;
assign addr[46599]= 1859775393;
assign addr[46600]= 1896833245;
assign addr[46601]= 1931484818;
assign addr[46602]= 1963686155;
assign addr[46603]= 1993396407;
assign addr[46604]= 2020577882;
assign addr[46605]= 2045196100;
assign addr[46606]= 2067219829;
assign addr[46607]= 2086621133;
assign addr[46608]= 2103375398;
assign addr[46609]= 2117461370;
assign addr[46610]= 2128861181;
assign addr[46611]= 2137560369;
assign addr[46612]= 2143547897;
assign addr[46613]= 2146816171;
assign addr[46614]= 2147361045;
assign addr[46615]= 2145181827;
assign addr[46616]= 2140281282;
assign addr[46617]= 2132665626;
assign addr[46618]= 2122344521;
assign addr[46619]= 2109331059;
assign addr[46620]= 2093641749;
assign addr[46621]= 2075296495;
assign addr[46622]= 2054318569;
assign addr[46623]= 2030734582;
assign addr[46624]= 2004574453;
assign addr[46625]= 1975871368;
assign addr[46626]= 1944661739;
assign addr[46627]= 1910985158;
assign addr[46628]= 1874884346;
assign addr[46629]= 1836405100;
assign addr[46630]= 1795596234;
assign addr[46631]= 1752509516;
assign addr[46632]= 1707199606;
assign addr[46633]= 1659723983;
assign addr[46634]= 1610142873;
assign addr[46635]= 1558519173;
assign addr[46636]= 1504918373;
assign addr[46637]= 1449408469;
assign addr[46638]= 1392059879;
assign addr[46639]= 1332945355;
assign addr[46640]= 1272139887;
assign addr[46641]= 1209720613;
assign addr[46642]= 1145766716;
assign addr[46643]= 1080359326;
assign addr[46644]= 1013581418;
assign addr[46645]= 945517704;
assign addr[46646]= 876254528;
assign addr[46647]= 805879757;
assign addr[46648]= 734482665;
assign addr[46649]= 662153826;
assign addr[46650]= 588984994;
assign addr[46651]= 515068990;
assign addr[46652]= 440499581;
assign addr[46653]= 365371365;
assign addr[46654]= 289779648;
assign addr[46655]= 213820322;
assign addr[46656]= 137589750;
assign addr[46657]= 61184634;
assign addr[46658]= -15298099;
assign addr[46659]= -91761426;
assign addr[46660]= -168108346;
assign addr[46661]= -244242007;
assign addr[46662]= -320065829;
assign addr[46663]= -395483624;
assign addr[46664]= -470399716;
assign addr[46665]= -544719071;
assign addr[46666]= -618347408;
assign addr[46667]= -691191324;
assign addr[46668]= -763158411;
assign addr[46669]= -834157373;
assign addr[46670]= -904098143;
assign addr[46671]= -972891995;
assign addr[46672]= -1040451659;
assign addr[46673]= -1106691431;
assign addr[46674]= -1171527280;
assign addr[46675]= -1234876957;
assign addr[46676]= -1296660098;
assign addr[46677]= -1356798326;
assign addr[46678]= -1415215352;
assign addr[46679]= -1471837070;
assign addr[46680]= -1526591649;
assign addr[46681]= -1579409630;
assign addr[46682]= -1630224009;
assign addr[46683]= -1678970324;
assign addr[46684]= -1725586737;
assign addr[46685]= -1770014111;
assign addr[46686]= -1812196087;
assign addr[46687]= -1852079154;
assign addr[46688]= -1889612716;
assign addr[46689]= -1924749160;
assign addr[46690]= -1957443913;
assign addr[46691]= -1987655498;
assign addr[46692]= -2015345591;
assign addr[46693]= -2040479063;
assign addr[46694]= -2063024031;
assign addr[46695]= -2082951896;
assign addr[46696]= -2100237377;
assign addr[46697]= -2114858546;
assign addr[46698]= -2126796855;
assign addr[46699]= -2136037160;
assign addr[46700]= -2142567738;
assign addr[46701]= -2146380306;
assign addr[46702]= -2147470025;
assign addr[46703]= -2145835515;
assign addr[46704]= -2141478848;
assign addr[46705]= -2134405552;
assign addr[46706]= -2124624598;
assign addr[46707]= -2112148396;
assign addr[46708]= -2096992772;
assign addr[46709]= -2079176953;
assign addr[46710]= -2058723538;
assign addr[46711]= -2035658475;
assign addr[46712]= -2010011024;
assign addr[46713]= -1981813720;
assign addr[46714]= -1951102334;
assign addr[46715]= -1917915825;
assign addr[46716]= -1882296293;
assign addr[46717]= -1844288924;
assign addr[46718]= -1803941934;
assign addr[46719]= -1761306505;
assign addr[46720]= -1716436725;
assign addr[46721]= -1669389513;
assign addr[46722]= -1620224553;
assign addr[46723]= -1569004214;
assign addr[46724]= -1515793473;
assign addr[46725]= -1460659832;
assign addr[46726]= -1403673233;
assign addr[46727]= -1344905966;
assign addr[46728]= -1284432584;
assign addr[46729]= -1222329801;
assign addr[46730]= -1158676398;
assign addr[46731]= -1093553126;
assign addr[46732]= -1027042599;
assign addr[46733]= -959229189;
assign addr[46734]= -890198924;
assign addr[46735]= -820039373;
assign addr[46736]= -748839539;
assign addr[46737]= -676689746;
assign addr[46738]= -603681519;
assign addr[46739]= -529907477;
assign addr[46740]= -455461206;
assign addr[46741]= -380437148;
assign addr[46742]= -304930476;
assign addr[46743]= -229036977;
assign addr[46744]= -152852926;
assign addr[46745]= -76474970;
assign addr[46746]= 0;
assign addr[46747]= 76474970;
assign addr[46748]= 152852926;
assign addr[46749]= 229036977;
assign addr[46750]= 304930476;
assign addr[46751]= 380437148;
assign addr[46752]= 455461206;
assign addr[46753]= 529907477;
assign addr[46754]= 603681519;
assign addr[46755]= 676689746;
assign addr[46756]= 748839539;
assign addr[46757]= 820039373;
assign addr[46758]= 890198924;
assign addr[46759]= 959229189;
assign addr[46760]= 1027042599;
assign addr[46761]= 1093553126;
assign addr[46762]= 1158676398;
assign addr[46763]= 1222329801;
assign addr[46764]= 1284432584;
assign addr[46765]= 1344905966;
assign addr[46766]= 1403673233;
assign addr[46767]= 1460659832;
assign addr[46768]= 1515793473;
assign addr[46769]= 1569004214;
assign addr[46770]= 1620224553;
assign addr[46771]= 1669389513;
assign addr[46772]= 1716436725;
assign addr[46773]= 1761306505;
assign addr[46774]= 1803941934;
assign addr[46775]= 1844288924;
assign addr[46776]= 1882296293;
assign addr[46777]= 1917915825;
assign addr[46778]= 1951102334;
assign addr[46779]= 1981813720;
assign addr[46780]= 2010011024;
assign addr[46781]= 2035658475;
assign addr[46782]= 2058723538;
assign addr[46783]= 2079176953;
assign addr[46784]= 2096992772;
assign addr[46785]= 2112148396;
assign addr[46786]= 2124624598;
assign addr[46787]= 2134405552;
assign addr[46788]= 2141478848;
assign addr[46789]= 2145835515;
assign addr[46790]= 2147470025;
assign addr[46791]= 2146380306;
assign addr[46792]= 2142567738;
assign addr[46793]= 2136037160;
assign addr[46794]= 2126796855;
assign addr[46795]= 2114858546;
assign addr[46796]= 2100237377;
assign addr[46797]= 2082951896;
assign addr[46798]= 2063024031;
assign addr[46799]= 2040479063;
assign addr[46800]= 2015345591;
assign addr[46801]= 1987655498;
assign addr[46802]= 1957443913;
assign addr[46803]= 1924749160;
assign addr[46804]= 1889612716;
assign addr[46805]= 1852079154;
assign addr[46806]= 1812196087;
assign addr[46807]= 1770014111;
assign addr[46808]= 1725586737;
assign addr[46809]= 1678970324;
assign addr[46810]= 1630224009;
assign addr[46811]= 1579409630;
assign addr[46812]= 1526591649;
assign addr[46813]= 1471837070;
assign addr[46814]= 1415215352;
assign addr[46815]= 1356798326;
assign addr[46816]= 1296660098;
assign addr[46817]= 1234876957;
assign addr[46818]= 1171527280;
assign addr[46819]= 1106691431;
assign addr[46820]= 1040451659;
assign addr[46821]= 972891995;
assign addr[46822]= 904098143;
assign addr[46823]= 834157373;
assign addr[46824]= 763158411;
assign addr[46825]= 691191324;
assign addr[46826]= 618347408;
assign addr[46827]= 544719071;
assign addr[46828]= 470399716;
assign addr[46829]= 395483624;
assign addr[46830]= 320065829;
assign addr[46831]= 244242007;
assign addr[46832]= 168108346;
assign addr[46833]= 91761426;
assign addr[46834]= 15298099;
assign addr[46835]= -61184634;
assign addr[46836]= -137589750;
assign addr[46837]= -213820322;
assign addr[46838]= -289779648;
assign addr[46839]= -365371365;
assign addr[46840]= -440499581;
assign addr[46841]= -515068990;
assign addr[46842]= -588984994;
assign addr[46843]= -662153826;
assign addr[46844]= -734482665;
assign addr[46845]= -805879757;
assign addr[46846]= -876254528;
assign addr[46847]= -945517704;
assign addr[46848]= -1013581418;
assign addr[46849]= -1080359326;
assign addr[46850]= -1145766716;
assign addr[46851]= -1209720613;
assign addr[46852]= -1272139887;
assign addr[46853]= -1332945355;
assign addr[46854]= -1392059879;
assign addr[46855]= -1449408469;
assign addr[46856]= -1504918373;
assign addr[46857]= -1558519173;
assign addr[46858]= -1610142873;
assign addr[46859]= -1659723983;
assign addr[46860]= -1707199606;
assign addr[46861]= -1752509516;
assign addr[46862]= -1795596234;
assign addr[46863]= -1836405100;
assign addr[46864]= -1874884346;
assign addr[46865]= -1910985158;
assign addr[46866]= -1944661739;
assign addr[46867]= -1975871368;
assign addr[46868]= -2004574453;
assign addr[46869]= -2030734582;
assign addr[46870]= -2054318569;
assign addr[46871]= -2075296495;
assign addr[46872]= -2093641749;
assign addr[46873]= -2109331059;
assign addr[46874]= -2122344521;
assign addr[46875]= -2132665626;
assign addr[46876]= -2140281282;
assign addr[46877]= -2145181827;
assign addr[46878]= -2147361045;
assign addr[46879]= -2146816171;
assign addr[46880]= -2143547897;
assign addr[46881]= -2137560369;
assign addr[46882]= -2128861181;
assign addr[46883]= -2117461370;
assign addr[46884]= -2103375398;
assign addr[46885]= -2086621133;
assign addr[46886]= -2067219829;
assign addr[46887]= -2045196100;
assign addr[46888]= -2020577882;
assign addr[46889]= -1993396407;
assign addr[46890]= -1963686155;
assign addr[46891]= -1931484818;
assign addr[46892]= -1896833245;
assign addr[46893]= -1859775393;
assign addr[46894]= -1820358275;
assign addr[46895]= -1778631892;
assign addr[46896]= -1734649179;
assign addr[46897]= -1688465931;
assign addr[46898]= -1640140734;
assign addr[46899]= -1589734894;
assign addr[46900]= -1537312353;
assign addr[46901]= -1482939614;
assign addr[46902]= -1426685652;
assign addr[46903]= -1368621831;
assign addr[46904]= -1308821808;
assign addr[46905]= -1247361445;
assign addr[46906]= -1184318708;
assign addr[46907]= -1119773573;
assign addr[46908]= -1053807919;
assign addr[46909]= -986505429;
assign addr[46910]= -917951481;
assign addr[46911]= -848233042;
assign addr[46912]= -777438554;
assign addr[46913]= -705657826;
assign addr[46914]= -632981917;
assign addr[46915]= -559503022;
assign addr[46916]= -485314355;
assign addr[46917]= -410510029;
assign addr[46918]= -335184940;
assign addr[46919]= -259434643;
assign addr[46920]= -183355234;
assign addr[46921]= -107043224;
assign addr[46922]= -30595422;
assign addr[46923]= 45891193;
assign addr[46924]= 122319591;
assign addr[46925]= 198592817;
assign addr[46926]= 274614114;
assign addr[46927]= 350287041;
assign addr[46928]= 425515602;
assign addr[46929]= 500204365;
assign addr[46930]= 574258580;
assign addr[46931]= 647584304;
assign addr[46932]= 720088517;
assign addr[46933]= 791679244;
assign addr[46934]= 862265664;
assign addr[46935]= 931758235;
assign addr[46936]= 1000068799;
assign addr[46937]= 1067110699;
assign addr[46938]= 1132798888;
assign addr[46939]= 1197050035;
assign addr[46940]= 1259782632;
assign addr[46941]= 1320917099;
assign addr[46942]= 1380375881;
assign addr[46943]= 1438083551;
assign addr[46944]= 1493966902;
assign addr[46945]= 1547955041;
assign addr[46946]= 1599979481;
assign addr[46947]= 1649974225;
assign addr[46948]= 1697875851;
assign addr[46949]= 1743623590;
assign addr[46950]= 1787159411;
assign addr[46951]= 1828428082;
assign addr[46952]= 1867377253;
assign addr[46953]= 1903957513;
assign addr[46954]= 1938122457;
assign addr[46955]= 1969828744;
assign addr[46956]= 1999036154;
assign addr[46957]= 2025707632;
assign addr[46958]= 2049809346;
assign addr[46959]= 2071310720;
assign addr[46960]= 2090184478;
assign addr[46961]= 2106406677;
assign addr[46962]= 2119956737;
assign addr[46963]= 2130817471;
assign addr[46964]= 2138975100;
assign addr[46965]= 2144419275;
assign addr[46966]= 2147143090;
assign addr[46967]= 2147143090;
assign addr[46968]= 2144419275;
assign addr[46969]= 2138975100;
assign addr[46970]= 2130817471;
assign addr[46971]= 2119956737;
assign addr[46972]= 2106406677;
assign addr[46973]= 2090184478;
assign addr[46974]= 2071310720;
assign addr[46975]= 2049809346;
assign addr[46976]= 2025707632;
assign addr[46977]= 1999036154;
assign addr[46978]= 1969828744;
assign addr[46979]= 1938122457;
assign addr[46980]= 1903957513;
assign addr[46981]= 1867377253;
assign addr[46982]= 1828428082;
assign addr[46983]= 1787159411;
assign addr[46984]= 1743623590;
assign addr[46985]= 1697875851;
assign addr[46986]= 1649974225;
assign addr[46987]= 1599979481;
assign addr[46988]= 1547955041;
assign addr[46989]= 1493966902;
assign addr[46990]= 1438083551;
assign addr[46991]= 1380375881;
assign addr[46992]= 1320917099;
assign addr[46993]= 1259782632;
assign addr[46994]= 1197050035;
assign addr[46995]= 1132798888;
assign addr[46996]= 1067110699;
assign addr[46997]= 1000068799;
assign addr[46998]= 931758235;
assign addr[46999]= 862265664;
assign addr[47000]= 791679244;
assign addr[47001]= 720088517;
assign addr[47002]= 647584304;
assign addr[47003]= 574258580;
assign addr[47004]= 500204365;
assign addr[47005]= 425515602;
assign addr[47006]= 350287041;
assign addr[47007]= 274614114;
assign addr[47008]= 198592817;
assign addr[47009]= 122319591;
assign addr[47010]= 45891193;
assign addr[47011]= -30595422;
assign addr[47012]= -107043224;
assign addr[47013]= -183355234;
assign addr[47014]= -259434643;
assign addr[47015]= -335184940;
assign addr[47016]= -410510029;
assign addr[47017]= -485314355;
assign addr[47018]= -559503022;
assign addr[47019]= -632981917;
assign addr[47020]= -705657826;
assign addr[47021]= -777438554;
assign addr[47022]= -848233042;
assign addr[47023]= -917951481;
assign addr[47024]= -986505429;
assign addr[47025]= -1053807919;
assign addr[47026]= -1119773573;
assign addr[47027]= -1184318708;
assign addr[47028]= -1247361445;
assign addr[47029]= -1308821808;
assign addr[47030]= -1368621831;
assign addr[47031]= -1426685652;
assign addr[47032]= -1482939614;
assign addr[47033]= -1537312353;
assign addr[47034]= -1589734894;
assign addr[47035]= -1640140734;
assign addr[47036]= -1688465931;
assign addr[47037]= -1734649179;
assign addr[47038]= -1778631892;
assign addr[47039]= -1820358275;
assign addr[47040]= -1859775393;
assign addr[47041]= -1896833245;
assign addr[47042]= -1931484818;
assign addr[47043]= -1963686155;
assign addr[47044]= -1993396407;
assign addr[47045]= -2020577882;
assign addr[47046]= -2045196100;
assign addr[47047]= -2067219829;
assign addr[47048]= -2086621133;
assign addr[47049]= -2103375398;
assign addr[47050]= -2117461370;
assign addr[47051]= -2128861181;
assign addr[47052]= -2137560369;
assign addr[47053]= -2143547897;
assign addr[47054]= -2146816171;
assign addr[47055]= -2147361045;
assign addr[47056]= -2145181827;
assign addr[47057]= -2140281282;
assign addr[47058]= -2132665626;
assign addr[47059]= -2122344521;
assign addr[47060]= -2109331059;
assign addr[47061]= -2093641749;
assign addr[47062]= -2075296495;
assign addr[47063]= -2054318569;
assign addr[47064]= -2030734582;
assign addr[47065]= -2004574453;
assign addr[47066]= -1975871368;
assign addr[47067]= -1944661739;
assign addr[47068]= -1910985158;
assign addr[47069]= -1874884346;
assign addr[47070]= -1836405100;
assign addr[47071]= -1795596234;
assign addr[47072]= -1752509516;
assign addr[47073]= -1707199606;
assign addr[47074]= -1659723983;
assign addr[47075]= -1610142873;
assign addr[47076]= -1558519173;
assign addr[47077]= -1504918373;
assign addr[47078]= -1449408469;
assign addr[47079]= -1392059879;
assign addr[47080]= -1332945355;
assign addr[47081]= -1272139887;
assign addr[47082]= -1209720613;
assign addr[47083]= -1145766716;
assign addr[47084]= -1080359326;
assign addr[47085]= -1013581418;
assign addr[47086]= -945517704;
assign addr[47087]= -876254528;
assign addr[47088]= -805879757;
assign addr[47089]= -734482665;
assign addr[47090]= -662153826;
assign addr[47091]= -588984994;
assign addr[47092]= -515068990;
assign addr[47093]= -440499581;
assign addr[47094]= -365371365;
assign addr[47095]= -289779648;
assign addr[47096]= -213820322;
assign addr[47097]= -137589750;
assign addr[47098]= -61184634;
assign addr[47099]= 15298099;
assign addr[47100]= 91761426;
assign addr[47101]= 168108346;
assign addr[47102]= 244242007;
assign addr[47103]= 320065829;
assign addr[47104]= 395483624;
assign addr[47105]= 470399716;
assign addr[47106]= 544719071;
assign addr[47107]= 618347408;
assign addr[47108]= 691191324;
assign addr[47109]= 763158411;
assign addr[47110]= 834157373;
assign addr[47111]= 904098143;
assign addr[47112]= 972891995;
assign addr[47113]= 1040451659;
assign addr[47114]= 1106691431;
assign addr[47115]= 1171527280;
assign addr[47116]= 1234876957;
assign addr[47117]= 1296660098;
assign addr[47118]= 1356798326;
assign addr[47119]= 1415215352;
assign addr[47120]= 1471837070;
assign addr[47121]= 1526591649;
assign addr[47122]= 1579409630;
assign addr[47123]= 1630224009;
assign addr[47124]= 1678970324;
assign addr[47125]= 1725586737;
assign addr[47126]= 1770014111;
assign addr[47127]= 1812196087;
assign addr[47128]= 1852079154;
assign addr[47129]= 1889612716;
assign addr[47130]= 1924749160;
assign addr[47131]= 1957443913;
assign addr[47132]= 1987655498;
assign addr[47133]= 2015345591;
assign addr[47134]= 2040479063;
assign addr[47135]= 2063024031;
assign addr[47136]= 2082951896;
assign addr[47137]= 2100237377;
assign addr[47138]= 2114858546;
assign addr[47139]= 2126796855;
assign addr[47140]= 2136037160;
assign addr[47141]= 2142567738;
assign addr[47142]= 2146380306;
assign addr[47143]= 2147470025;
assign addr[47144]= 2145835515;
assign addr[47145]= 2141478848;
assign addr[47146]= 2134405552;
assign addr[47147]= 2124624598;
assign addr[47148]= 2112148396;
assign addr[47149]= 2096992772;
assign addr[47150]= 2079176953;
assign addr[47151]= 2058723538;
assign addr[47152]= 2035658475;
assign addr[47153]= 2010011024;
assign addr[47154]= 1981813720;
assign addr[47155]= 1951102334;
assign addr[47156]= 1917915825;
assign addr[47157]= 1882296293;
assign addr[47158]= 1844288924;
assign addr[47159]= 1803941934;
assign addr[47160]= 1761306505;
assign addr[47161]= 1716436725;
assign addr[47162]= 1669389513;
assign addr[47163]= 1620224553;
assign addr[47164]= 1569004214;
assign addr[47165]= 1515793473;
assign addr[47166]= 1460659832;
assign addr[47167]= 1403673233;
assign addr[47168]= 1344905966;
assign addr[47169]= 1284432584;
assign addr[47170]= 1222329801;
assign addr[47171]= 1158676398;
assign addr[47172]= 1093553126;
assign addr[47173]= 1027042599;
assign addr[47174]= 959229189;
assign addr[47175]= 890198924;
assign addr[47176]= 820039373;
assign addr[47177]= 748839539;
assign addr[47178]= 676689746;
assign addr[47179]= 603681519;
assign addr[47180]= 529907477;
assign addr[47181]= 455461206;
assign addr[47182]= 380437148;
assign addr[47183]= 304930476;
assign addr[47184]= 229036977;
assign addr[47185]= 152852926;
assign addr[47186]= 76474970;
assign addr[47187]= 0;
assign addr[47188]= -76474970;
assign addr[47189]= -152852926;
assign addr[47190]= -229036977;
assign addr[47191]= -304930476;
assign addr[47192]= -380437148;
assign addr[47193]= -455461206;
assign addr[47194]= -529907477;
assign addr[47195]= -603681519;
assign addr[47196]= -676689746;
assign addr[47197]= -748839539;
assign addr[47198]= -820039373;
assign addr[47199]= -890198924;
assign addr[47200]= -959229189;
assign addr[47201]= -1027042599;
assign addr[47202]= -1093553126;
assign addr[47203]= -1158676398;
assign addr[47204]= -1222329801;
assign addr[47205]= -1284432584;
assign addr[47206]= -1344905966;
assign addr[47207]= -1403673233;
assign addr[47208]= -1460659832;
assign addr[47209]= -1515793473;
assign addr[47210]= -1569004214;
assign addr[47211]= -1620224553;
assign addr[47212]= -1669389513;
assign addr[47213]= -1716436725;
assign addr[47214]= -1761306505;
assign addr[47215]= -1803941934;
assign addr[47216]= -1844288924;
assign addr[47217]= -1882296293;
assign addr[47218]= -1917915825;
assign addr[47219]= -1951102334;
assign addr[47220]= -1981813720;
assign addr[47221]= -2010011024;
assign addr[47222]= -2035658475;
assign addr[47223]= -2058723538;
assign addr[47224]= -2079176953;
assign addr[47225]= -2096992772;
assign addr[47226]= -2112148396;
assign addr[47227]= -2124624598;
assign addr[47228]= -2134405552;
assign addr[47229]= -2141478848;
assign addr[47230]= -2145835515;
assign addr[47231]= -2147470025;
assign addr[47232]= -2146380306;
assign addr[47233]= -2142567738;
assign addr[47234]= -2136037160;
assign addr[47235]= -2126796855;
assign addr[47236]= -2114858546;
assign addr[47237]= -2100237377;
assign addr[47238]= -2082951896;
assign addr[47239]= -2063024031;
assign addr[47240]= -2040479063;
assign addr[47241]= -2015345591;
assign addr[47242]= -1987655498;
assign addr[47243]= -1957443913;
assign addr[47244]= -1924749160;
assign addr[47245]= -1889612716;
assign addr[47246]= -1852079154;
assign addr[47247]= -1812196087;
assign addr[47248]= -1770014111;
assign addr[47249]= -1725586737;
assign addr[47250]= -1678970324;
assign addr[47251]= -1630224009;
assign addr[47252]= -1579409630;
assign addr[47253]= -1526591649;
assign addr[47254]= -1471837070;
assign addr[47255]= -1415215352;
assign addr[47256]= -1356798326;
assign addr[47257]= -1296660098;
assign addr[47258]= -1234876957;
assign addr[47259]= -1171527280;
assign addr[47260]= -1106691431;
assign addr[47261]= -1040451659;
assign addr[47262]= -972891995;
assign addr[47263]= -904098143;
assign addr[47264]= -834157373;
assign addr[47265]= -763158411;
assign addr[47266]= -691191324;
assign addr[47267]= -618347408;
assign addr[47268]= -544719071;
assign addr[47269]= -470399716;
assign addr[47270]= -395483624;
assign addr[47271]= -320065829;
assign addr[47272]= -244242007;
assign addr[47273]= -168108346;
assign addr[47274]= -91761426;
assign addr[47275]= -15298099;
assign addr[47276]= 61184634;
assign addr[47277]= 137589750;
assign addr[47278]= 213820322;
assign addr[47279]= 289779648;
assign addr[47280]= 365371365;
assign addr[47281]= 440499581;
assign addr[47282]= 515068990;
assign addr[47283]= 588984994;
assign addr[47284]= 662153826;
assign addr[47285]= 734482665;
assign addr[47286]= 805879757;
assign addr[47287]= 876254528;
assign addr[47288]= 945517704;
assign addr[47289]= 1013581418;
assign addr[47290]= 1080359326;
assign addr[47291]= 1145766716;
assign addr[47292]= 1209720613;
assign addr[47293]= 1272139887;
assign addr[47294]= 1332945355;
assign addr[47295]= 1392059879;
assign addr[47296]= 1449408469;
assign addr[47297]= 1504918373;
assign addr[47298]= 1558519173;
assign addr[47299]= 1610142873;
assign addr[47300]= 1659723983;
assign addr[47301]= 1707199606;
assign addr[47302]= 1752509516;
assign addr[47303]= 1795596234;
assign addr[47304]= 1836405100;
assign addr[47305]= 1874884346;
assign addr[47306]= 1910985158;
assign addr[47307]= 1944661739;
assign addr[47308]= 1975871368;
assign addr[47309]= 2004574453;
assign addr[47310]= 2030734582;
assign addr[47311]= 2054318569;
assign addr[47312]= 2075296495;
assign addr[47313]= 2093641749;
assign addr[47314]= 2109331059;
assign addr[47315]= 2122344521;
assign addr[47316]= 2132665626;
assign addr[47317]= 2140281282;
assign addr[47318]= 2145181827;
assign addr[47319]= 2147361045;
assign addr[47320]= 2146816171;
assign addr[47321]= 2143547897;
assign addr[47322]= 2137560369;
assign addr[47323]= 2128861181;
assign addr[47324]= 2117461370;
assign addr[47325]= 2103375398;
assign addr[47326]= 2086621133;
assign addr[47327]= 2067219829;
assign addr[47328]= 2045196100;
assign addr[47329]= 2020577882;
assign addr[47330]= 1993396407;
assign addr[47331]= 1963686155;
assign addr[47332]= 1931484818;
assign addr[47333]= 1896833245;
assign addr[47334]= 1859775393;
assign addr[47335]= 1820358275;
assign addr[47336]= 1778631892;
assign addr[47337]= 1734649179;
assign addr[47338]= 1688465931;
assign addr[47339]= 1640140734;
assign addr[47340]= 1589734894;
assign addr[47341]= 1537312353;
assign addr[47342]= 1482939614;
assign addr[47343]= 1426685652;
assign addr[47344]= 1368621831;
assign addr[47345]= 1308821808;
assign addr[47346]= 1247361445;
assign addr[47347]= 1184318708;
assign addr[47348]= 1119773573;
assign addr[47349]= 1053807919;
assign addr[47350]= 986505429;
assign addr[47351]= 917951481;
assign addr[47352]= 848233042;
assign addr[47353]= 777438554;
assign addr[47354]= 705657826;
assign addr[47355]= 632981917;
assign addr[47356]= 559503022;
assign addr[47357]= 485314355;
assign addr[47358]= 410510029;
assign addr[47359]= 335184940;
assign addr[47360]= 259434643;
assign addr[47361]= 183355234;
assign addr[47362]= 107043224;
assign addr[47363]= 30595422;
assign addr[47364]= -45891193;
assign addr[47365]= -122319591;
assign addr[47366]= -198592817;
assign addr[47367]= -274614114;
assign addr[47368]= -350287041;
assign addr[47369]= -425515602;
assign addr[47370]= -500204365;
assign addr[47371]= -574258580;
assign addr[47372]= -647584304;
assign addr[47373]= -720088517;
assign addr[47374]= -791679244;
assign addr[47375]= -862265664;
assign addr[47376]= -931758235;
assign addr[47377]= -1000068799;
assign addr[47378]= -1067110699;
assign addr[47379]= -1132798888;
assign addr[47380]= -1197050035;
assign addr[47381]= -1259782632;
assign addr[47382]= -1320917099;
assign addr[47383]= -1380375881;
assign addr[47384]= -1438083551;
assign addr[47385]= -1493966902;
assign addr[47386]= -1547955041;
assign addr[47387]= -1599979481;
assign addr[47388]= -1649974225;
assign addr[47389]= -1697875851;
assign addr[47390]= -1743623590;
assign addr[47391]= -1787159411;
assign addr[47392]= -1828428082;
assign addr[47393]= -1867377253;
assign addr[47394]= -1903957513;
assign addr[47395]= -1938122457;
assign addr[47396]= -1969828744;
assign addr[47397]= -1999036154;
assign addr[47398]= -2025707632;
assign addr[47399]= -2049809346;
assign addr[47400]= -2071310720;
assign addr[47401]= -2090184478;
assign addr[47402]= -2106406677;
assign addr[47403]= -2119956737;
assign addr[47404]= -2130817471;
assign addr[47405]= -2138975100;
assign addr[47406]= -2144419275;
assign addr[47407]= -2147143090;
assign addr[47408]= -2147143090;
assign addr[47409]= -2144419275;
assign addr[47410]= -2138975100;
assign addr[47411]= -2130817471;
assign addr[47412]= -2119956737;
assign addr[47413]= -2106406677;
assign addr[47414]= -2090184478;
assign addr[47415]= -2071310720;
assign addr[47416]= -2049809346;
assign addr[47417]= -2025707632;
assign addr[47418]= -1999036154;
assign addr[47419]= -1969828744;
assign addr[47420]= -1938122457;
assign addr[47421]= -1903957513;
assign addr[47422]= -1867377253;
assign addr[47423]= -1828428082;
assign addr[47424]= -1787159411;
assign addr[47425]= -1743623590;
assign addr[47426]= -1697875851;
assign addr[47427]= -1649974225;
assign addr[47428]= -1599979481;
assign addr[47429]= -1547955041;
assign addr[47430]= -1493966902;
assign addr[47431]= -1438083551;
assign addr[47432]= -1380375881;
assign addr[47433]= -1320917099;
assign addr[47434]= -1259782632;
assign addr[47435]= -1197050035;
assign addr[47436]= -1132798888;
assign addr[47437]= -1067110699;
assign addr[47438]= -1000068799;
assign addr[47439]= -931758235;
assign addr[47440]= -862265664;
assign addr[47441]= -791679244;
assign addr[47442]= -720088517;
assign addr[47443]= -647584304;
assign addr[47444]= -574258580;
assign addr[47445]= -500204365;
assign addr[47446]= -425515602;
assign addr[47447]= -350287041;
assign addr[47448]= -274614114;
assign addr[47449]= -198592817;
assign addr[47450]= -122319591;
assign addr[47451]= -45891193;
assign addr[47452]= 30595422;
assign addr[47453]= 107043224;
assign addr[47454]= 183355234;
assign addr[47455]= 259434643;
assign addr[47456]= 335184940;
assign addr[47457]= 410510029;
assign addr[47458]= 485314355;
assign addr[47459]= 559503022;
assign addr[47460]= 632981917;
assign addr[47461]= 705657826;
assign addr[47462]= 777438554;
assign addr[47463]= 848233042;
assign addr[47464]= 917951481;
assign addr[47465]= 986505429;
assign addr[47466]= 1053807919;
assign addr[47467]= 1119773573;
assign addr[47468]= 1184318708;
assign addr[47469]= 1247361445;
assign addr[47470]= 1308821808;
assign addr[47471]= 1368621831;
assign addr[47472]= 1426685652;
assign addr[47473]= 1482939614;
assign addr[47474]= 1537312353;
assign addr[47475]= 1589734894;
assign addr[47476]= 1640140734;
assign addr[47477]= 1688465931;
assign addr[47478]= 1734649179;
assign addr[47479]= 1778631892;
assign addr[47480]= 1820358275;
assign addr[47481]= 1859775393;
assign addr[47482]= 1896833245;
assign addr[47483]= 1931484818;
assign addr[47484]= 1963686155;
assign addr[47485]= 1993396407;
assign addr[47486]= 2020577882;
assign addr[47487]= 2045196100;
assign addr[47488]= 2067219829;
assign addr[47489]= 2086621133;
assign addr[47490]= 2103375398;
assign addr[47491]= 2117461370;
assign addr[47492]= 2128861181;
assign addr[47493]= 2137560369;
assign addr[47494]= 2143547897;
assign addr[47495]= 2146816171;
assign addr[47496]= 2147361045;
assign addr[47497]= 2145181827;
assign addr[47498]= 2140281282;
assign addr[47499]= 2132665626;
assign addr[47500]= 2122344521;
assign addr[47501]= 2109331059;
assign addr[47502]= 2093641749;
assign addr[47503]= 2075296495;
assign addr[47504]= 2054318569;
assign addr[47505]= 2030734582;
assign addr[47506]= 2004574453;
assign addr[47507]= 1975871368;
assign addr[47508]= 1944661739;
assign addr[47509]= 1910985158;
assign addr[47510]= 1874884346;
assign addr[47511]= 1836405100;
assign addr[47512]= 1795596234;
assign addr[47513]= 1752509516;
assign addr[47514]= 1707199606;
assign addr[47515]= 1659723983;
assign addr[47516]= 1610142873;
assign addr[47517]= 1558519173;
assign addr[47518]= 1504918373;
assign addr[47519]= 1449408469;
assign addr[47520]= 1392059879;
assign addr[47521]= 1332945355;
assign addr[47522]= 1272139887;
assign addr[47523]= 1209720613;
assign addr[47524]= 1145766716;
assign addr[47525]= 1080359326;
assign addr[47526]= 1013581418;
assign addr[47527]= 945517704;
assign addr[47528]= 876254528;
assign addr[47529]= 805879757;
assign addr[47530]= 734482665;
assign addr[47531]= 662153826;
assign addr[47532]= 588984994;
assign addr[47533]= 515068990;
assign addr[47534]= 440499581;
assign addr[47535]= 365371365;
assign addr[47536]= 289779648;
assign addr[47537]= 213820322;
assign addr[47538]= 137589750;
assign addr[47539]= 61184634;
assign addr[47540]= -15298099;
assign addr[47541]= -91761426;
assign addr[47542]= -168108346;
assign addr[47543]= -244242007;
assign addr[47544]= -320065829;
assign addr[47545]= -395483624;
assign addr[47546]= -470399716;
assign addr[47547]= -544719071;
assign addr[47548]= -618347408;
assign addr[47549]= -691191324;
assign addr[47550]= -763158411;
assign addr[47551]= -834157373;
assign addr[47552]= -904098143;
assign addr[47553]= -972891995;
assign addr[47554]= -1040451659;
assign addr[47555]= -1106691431;
assign addr[47556]= -1171527280;
assign addr[47557]= -1234876957;
assign addr[47558]= -1296660098;
assign addr[47559]= -1356798326;
assign addr[47560]= -1415215352;
assign addr[47561]= -1471837070;
assign addr[47562]= -1526591649;
assign addr[47563]= -1579409630;
assign addr[47564]= -1630224009;
assign addr[47565]= -1678970324;
assign addr[47566]= -1725586737;
assign addr[47567]= -1770014111;
assign addr[47568]= -1812196087;
assign addr[47569]= -1852079154;
assign addr[47570]= -1889612716;
assign addr[47571]= -1924749160;
assign addr[47572]= -1957443913;
assign addr[47573]= -1987655498;
assign addr[47574]= -2015345591;
assign addr[47575]= -2040479063;
assign addr[47576]= -2063024031;
assign addr[47577]= -2082951896;
assign addr[47578]= -2100237377;
assign addr[47579]= -2114858546;
assign addr[47580]= -2126796855;
assign addr[47581]= -2136037160;
assign addr[47582]= -2142567738;
assign addr[47583]= -2146380306;
assign addr[47584]= -2147470025;
assign addr[47585]= -2145835515;
assign addr[47586]= -2141478848;
assign addr[47587]= -2134405552;
assign addr[47588]= -2124624598;
assign addr[47589]= -2112148396;
assign addr[47590]= -2096992772;
assign addr[47591]= -2079176953;
assign addr[47592]= -2058723538;
assign addr[47593]= -2035658475;
assign addr[47594]= -2010011024;
assign addr[47595]= -1981813720;
assign addr[47596]= -1951102334;
assign addr[47597]= -1917915825;
assign addr[47598]= -1882296293;
assign addr[47599]= -1844288924;
assign addr[47600]= -1803941934;
assign addr[47601]= -1761306505;
assign addr[47602]= -1716436725;
assign addr[47603]= -1669389513;
assign addr[47604]= -1620224553;
assign addr[47605]= -1569004214;
assign addr[47606]= -1515793473;
assign addr[47607]= -1460659832;
assign addr[47608]= -1403673233;
assign addr[47609]= -1344905966;
assign addr[47610]= -1284432584;
assign addr[47611]= -1222329801;
assign addr[47612]= -1158676398;
assign addr[47613]= -1093553126;
assign addr[47614]= -1027042599;
assign addr[47615]= -959229189;
assign addr[47616]= -890198924;
assign addr[47617]= -820039373;
assign addr[47618]= -748839539;
assign addr[47619]= -676689746;
assign addr[47620]= -603681519;
assign addr[47621]= -529907477;
assign addr[47622]= -455461206;
assign addr[47623]= -380437148;
assign addr[47624]= -304930476;
assign addr[47625]= -229036977;
assign addr[47626]= -152852926;
assign addr[47627]= -76474970;
assign addr[47628]= 0;
assign addr[47629]= 76474970;
assign addr[47630]= 152852926;
assign addr[47631]= 229036977;
assign addr[47632]= 304930476;
assign addr[47633]= 380437148;
assign addr[47634]= 455461206;
assign addr[47635]= 529907477;
assign addr[47636]= 603681519;
assign addr[47637]= 676689746;
assign addr[47638]= 748839539;
assign addr[47639]= 820039373;
assign addr[47640]= 890198924;
assign addr[47641]= 959229189;
assign addr[47642]= 1027042599;
assign addr[47643]= 1093553126;
assign addr[47644]= 1158676398;
assign addr[47645]= 1222329801;
assign addr[47646]= 1284432584;
assign addr[47647]= 1344905966;
assign addr[47648]= 1403673233;
assign addr[47649]= 1460659832;
assign addr[47650]= 1515793473;
assign addr[47651]= 1569004214;
assign addr[47652]= 1620224553;
assign addr[47653]= 1669389513;
assign addr[47654]= 1716436725;
assign addr[47655]= 1761306505;
assign addr[47656]= 1803941934;
assign addr[47657]= 1844288924;
assign addr[47658]= 1882296293;
assign addr[47659]= 1917915825;
assign addr[47660]= 1951102334;
assign addr[47661]= 1981813720;
assign addr[47662]= 2010011024;
assign addr[47663]= 2035658475;
assign addr[47664]= 2058723538;
assign addr[47665]= 2079176953;
assign addr[47666]= 2096992772;
assign addr[47667]= 2112148396;
assign addr[47668]= 2124624598;
assign addr[47669]= 2134405552;
assign addr[47670]= 2141478848;
assign addr[47671]= 2145835515;
assign addr[47672]= 2147470025;
assign addr[47673]= 2146380306;
assign addr[47674]= 2142567738;
assign addr[47675]= 2136037160;
assign addr[47676]= 2126796855;
assign addr[47677]= 2114858546;
assign addr[47678]= 2100237377;
assign addr[47679]= 2082951896;
assign addr[47680]= 2063024031;
assign addr[47681]= 2040479063;
assign addr[47682]= 2015345591;
assign addr[47683]= 1987655498;
assign addr[47684]= 1957443913;
assign addr[47685]= 1924749160;
assign addr[47686]= 1889612716;
assign addr[47687]= 1852079154;
assign addr[47688]= 1812196087;
assign addr[47689]= 1770014111;
assign addr[47690]= 1725586737;
assign addr[47691]= 1678970324;
assign addr[47692]= 1630224009;
assign addr[47693]= 1579409630;
assign addr[47694]= 1526591649;
assign addr[47695]= 1471837070;
assign addr[47696]= 1415215352;
assign addr[47697]= 1356798326;
assign addr[47698]= 1296660098;
assign addr[47699]= 1234876957;
assign addr[47700]= 1171527280;
assign addr[47701]= 1106691431;
assign addr[47702]= 1040451659;
assign addr[47703]= 972891995;
assign addr[47704]= 904098143;
assign addr[47705]= 834157373;
assign addr[47706]= 763158411;
assign addr[47707]= 691191324;
assign addr[47708]= 618347408;
assign addr[47709]= 544719071;
assign addr[47710]= 470399716;
assign addr[47711]= 395483624;
assign addr[47712]= 320065829;
assign addr[47713]= 244242007;
assign addr[47714]= 168108346;
assign addr[47715]= 91761426;
assign addr[47716]= 15298099;
assign addr[47717]= -61184634;
assign addr[47718]= -137589750;
assign addr[47719]= -213820322;
assign addr[47720]= -289779648;
assign addr[47721]= -365371365;
assign addr[47722]= -440499581;
assign addr[47723]= -515068990;
assign addr[47724]= -588984994;
assign addr[47725]= -662153826;
assign addr[47726]= -734482665;
assign addr[47727]= -805879757;
assign addr[47728]= -876254528;
assign addr[47729]= -945517704;
assign addr[47730]= -1013581418;
assign addr[47731]= -1080359326;
assign addr[47732]= -1145766716;
assign addr[47733]= -1209720613;
assign addr[47734]= -1272139887;
assign addr[47735]= -1332945355;
assign addr[47736]= -1392059879;
assign addr[47737]= -1449408469;
assign addr[47738]= -1504918373;
assign addr[47739]= -1558519173;
assign addr[47740]= -1610142873;
assign addr[47741]= -1659723983;
assign addr[47742]= -1707199606;
assign addr[47743]= -1752509516;
assign addr[47744]= -1795596234;
assign addr[47745]= -1836405100;
assign addr[47746]= -1874884346;
assign addr[47747]= -1910985158;
assign addr[47748]= -1944661739;
assign addr[47749]= -1975871368;
assign addr[47750]= -2004574453;
assign addr[47751]= -2030734582;
assign addr[47752]= -2054318569;
assign addr[47753]= -2075296495;
assign addr[47754]= -2093641749;
assign addr[47755]= -2109331059;
assign addr[47756]= -2122344521;
assign addr[47757]= -2132665626;
assign addr[47758]= -2140281282;
assign addr[47759]= -2145181827;
assign addr[47760]= -2147361045;
assign addr[47761]= -2146816171;
assign addr[47762]= -2143547897;
assign addr[47763]= -2137560369;
assign addr[47764]= -2128861181;
assign addr[47765]= -2117461370;
assign addr[47766]= -2103375398;
assign addr[47767]= -2086621133;
assign addr[47768]= -2067219829;
assign addr[47769]= -2045196100;
assign addr[47770]= -2020577882;
assign addr[47771]= -1993396407;
assign addr[47772]= -1963686155;
assign addr[47773]= -1931484818;
assign addr[47774]= -1896833245;
assign addr[47775]= -1859775393;
assign addr[47776]= -1820358275;
assign addr[47777]= -1778631892;
assign addr[47778]= -1734649179;
assign addr[47779]= -1688465931;
assign addr[47780]= -1640140734;
assign addr[47781]= -1589734894;
assign addr[47782]= -1537312353;
assign addr[47783]= -1482939614;
assign addr[47784]= -1426685652;
assign addr[47785]= -1368621831;
assign addr[47786]= -1308821808;
assign addr[47787]= -1247361445;
assign addr[47788]= -1184318708;
assign addr[47789]= -1119773573;
assign addr[47790]= -1053807919;
assign addr[47791]= -986505429;
assign addr[47792]= -917951481;
assign addr[47793]= -848233042;
assign addr[47794]= -777438554;
assign addr[47795]= -705657826;
assign addr[47796]= -632981917;
assign addr[47797]= -559503022;
assign addr[47798]= -485314355;
assign addr[47799]= -410510029;
assign addr[47800]= -335184940;
assign addr[47801]= -259434643;
assign addr[47802]= -183355234;
assign addr[47803]= -107043224;
assign addr[47804]= -30595422;
assign addr[47805]= 45891193;
assign addr[47806]= 122319591;
assign addr[47807]= 198592817;
assign addr[47808]= 274614114;
assign addr[47809]= 350287041;
assign addr[47810]= 425515602;
assign addr[47811]= 500204365;
assign addr[47812]= 574258580;
assign addr[47813]= 647584304;
assign addr[47814]= 720088517;
assign addr[47815]= 791679244;
assign addr[47816]= 862265664;
assign addr[47817]= 931758235;
assign addr[47818]= 1000068799;
assign addr[47819]= 1067110699;
assign addr[47820]= 1132798888;
assign addr[47821]= 1197050035;
assign addr[47822]= 1259782632;
assign addr[47823]= 1320917099;
assign addr[47824]= 1380375881;
assign addr[47825]= 1438083551;
assign addr[47826]= 1493966902;
assign addr[47827]= 1547955041;
assign addr[47828]= 1599979481;
assign addr[47829]= 1649974225;
assign addr[47830]= 1697875851;
assign addr[47831]= 1743623590;
assign addr[47832]= 1787159411;
assign addr[47833]= 1828428082;
assign addr[47834]= 1867377253;
assign addr[47835]= 1903957513;
assign addr[47836]= 1938122457;
assign addr[47837]= 1969828744;
assign addr[47838]= 1999036154;
assign addr[47839]= 2025707632;
assign addr[47840]= 2049809346;
assign addr[47841]= 2071310720;
assign addr[47842]= 2090184478;
assign addr[47843]= 2106406677;
assign addr[47844]= 2119956737;
assign addr[47845]= 2130817471;
assign addr[47846]= 2138975100;
assign addr[47847]= 2144419275;
assign addr[47848]= 2147143090;
assign addr[47849]= 2147143090;
assign addr[47850]= 2144419275;
assign addr[47851]= 2138975100;
assign addr[47852]= 2130817471;
assign addr[47853]= 2119956737;
assign addr[47854]= 2106406677;
assign addr[47855]= 2090184478;
assign addr[47856]= 2071310720;
assign addr[47857]= 2049809346;
assign addr[47858]= 2025707632;
assign addr[47859]= 1999036154;
assign addr[47860]= 1969828744;
assign addr[47861]= 1938122457;
assign addr[47862]= 1903957513;
assign addr[47863]= 1867377253;
assign addr[47864]= 1828428082;
assign addr[47865]= 1787159411;
assign addr[47866]= 1743623590;
assign addr[47867]= 1697875851;
assign addr[47868]= 1649974225;
assign addr[47869]= 1599979481;
assign addr[47870]= 1547955041;
assign addr[47871]= 1493966902;
assign addr[47872]= 1438083551;
assign addr[47873]= 1380375881;
assign addr[47874]= 1320917099;
assign addr[47875]= 1259782632;
assign addr[47876]= 1197050035;
assign addr[47877]= 1132798888;
assign addr[47878]= 1067110699;
assign addr[47879]= 1000068799;
assign addr[47880]= 931758235;
assign addr[47881]= 862265664;
assign addr[47882]= 791679244;
assign addr[47883]= 720088517;
assign addr[47884]= 647584304;
assign addr[47885]= 574258580;
assign addr[47886]= 500204365;
assign addr[47887]= 425515602;
assign addr[47888]= 350287041;
assign addr[47889]= 274614114;
assign addr[47890]= 198592817;
assign addr[47891]= 122319591;
assign addr[47892]= 45891193;
assign addr[47893]= -30595422;
assign addr[47894]= -107043224;
assign addr[47895]= -183355234;
assign addr[47896]= -259434643;
assign addr[47897]= -335184940;
assign addr[47898]= -410510029;
assign addr[47899]= -485314355;
assign addr[47900]= -559503022;
assign addr[47901]= -632981917;
assign addr[47902]= -705657826;
assign addr[47903]= -777438554;
assign addr[47904]= -848233042;
assign addr[47905]= -917951481;
assign addr[47906]= -986505429;
assign addr[47907]= -1053807919;
assign addr[47908]= -1119773573;
assign addr[47909]= -1184318708;
assign addr[47910]= -1247361445;
assign addr[47911]= -1308821808;
assign addr[47912]= -1368621831;
assign addr[47913]= -1426685652;
assign addr[47914]= -1482939614;
assign addr[47915]= -1537312353;
assign addr[47916]= -1589734894;
assign addr[47917]= -1640140734;
assign addr[47918]= -1688465931;
assign addr[47919]= -1734649179;
assign addr[47920]= -1778631892;
assign addr[47921]= -1820358275;
assign addr[47922]= -1859775393;
assign addr[47923]= -1896833245;
assign addr[47924]= -1931484818;
assign addr[47925]= -1963686155;
assign addr[47926]= -1993396407;
assign addr[47927]= -2020577882;
assign addr[47928]= -2045196100;
assign addr[47929]= -2067219829;
assign addr[47930]= -2086621133;
assign addr[47931]= -2103375398;
assign addr[47932]= -2117461370;
assign addr[47933]= -2128861181;
assign addr[47934]= -2137560369;
assign addr[47935]= -2143547897;
assign addr[47936]= -2146816171;
assign addr[47937]= -2147361045;
assign addr[47938]= -2145181827;
assign addr[47939]= -2140281282;
assign addr[47940]= -2132665626;
assign addr[47941]= -2122344521;
assign addr[47942]= -2109331059;
assign addr[47943]= -2093641749;
assign addr[47944]= -2075296495;
assign addr[47945]= -2054318569;
assign addr[47946]= -2030734582;
assign addr[47947]= -2004574453;
assign addr[47948]= -1975871368;
assign addr[47949]= -1944661739;
assign addr[47950]= -1910985158;
assign addr[47951]= -1874884346;
assign addr[47952]= -1836405100;
assign addr[47953]= -1795596234;
assign addr[47954]= -1752509516;
assign addr[47955]= -1707199606;
assign addr[47956]= -1659723983;
assign addr[47957]= -1610142873;
assign addr[47958]= -1558519173;
assign addr[47959]= -1504918373;
assign addr[47960]= -1449408469;
assign addr[47961]= -1392059879;
assign addr[47962]= -1332945355;
assign addr[47963]= -1272139887;
assign addr[47964]= -1209720613;
assign addr[47965]= -1145766716;
assign addr[47966]= -1080359326;
assign addr[47967]= -1013581418;
assign addr[47968]= -945517704;
assign addr[47969]= -876254528;
assign addr[47970]= -805879757;
assign addr[47971]= -734482665;
assign addr[47972]= -662153826;
assign addr[47973]= -588984994;
assign addr[47974]= -515068990;
assign addr[47975]= -440499581;
assign addr[47976]= -365371365;
assign addr[47977]= -289779648;
assign addr[47978]= -213820322;
assign addr[47979]= -137589750;
assign addr[47980]= -61184634;
assign addr[47981]= 15298099;
assign addr[47982]= 91761426;
assign addr[47983]= 168108346;
assign addr[47984]= 244242007;
assign addr[47985]= 320065829;
assign addr[47986]= 395483624;
assign addr[47987]= 470399716;
assign addr[47988]= 544719071;
assign addr[47989]= 618347408;
assign addr[47990]= 691191324;
assign addr[47991]= 763158411;
assign addr[47992]= 834157373;
assign addr[47993]= 904098143;
assign addr[47994]= 972891995;
assign addr[47995]= 1040451659;
assign addr[47996]= 1106691431;
assign addr[47997]= 1171527280;
assign addr[47998]= 1234876957;
assign addr[47999]= 1296660098;
assign addr[48000]= 1356798326;
assign addr[48001]= 1415215352;
assign addr[48002]= 1471837070;
assign addr[48003]= 1526591649;
assign addr[48004]= 1579409630;
assign addr[48005]= 1630224009;
assign addr[48006]= 1678970324;
assign addr[48007]= 1725586737;
assign addr[48008]= 1770014111;
assign addr[48009]= 1812196087;
assign addr[48010]= 1852079154;
assign addr[48011]= 1889612716;
assign addr[48012]= 1924749160;
assign addr[48013]= 1957443913;
assign addr[48014]= 1987655498;
assign addr[48015]= 2015345591;
assign addr[48016]= 2040479063;
assign addr[48017]= 2063024031;
assign addr[48018]= 2082951896;
assign addr[48019]= 2100237377;
assign addr[48020]= 2114858546;
assign addr[48021]= 2126796855;
assign addr[48022]= 2136037160;
assign addr[48023]= 2142567738;
assign addr[48024]= 2146380306;
assign addr[48025]= 2147470025;
assign addr[48026]= 2145835515;
assign addr[48027]= 2141478848;
assign addr[48028]= 2134405552;
assign addr[48029]= 2124624598;
assign addr[48030]= 2112148396;
assign addr[48031]= 2096992772;
assign addr[48032]= 2079176953;
assign addr[48033]= 2058723538;
assign addr[48034]= 2035658475;
assign addr[48035]= 2010011024;
assign addr[48036]= 1981813720;
assign addr[48037]= 1951102334;
assign addr[48038]= 1917915825;
assign addr[48039]= 1882296293;
assign addr[48040]= 1844288924;
assign addr[48041]= 1803941934;
assign addr[48042]= 1761306505;
assign addr[48043]= 1716436725;
assign addr[48044]= 1669389513;
assign addr[48045]= 1620224553;
assign addr[48046]= 1569004214;
assign addr[48047]= 1515793473;
assign addr[48048]= 1460659832;
assign addr[48049]= 1403673233;
assign addr[48050]= 1344905966;
assign addr[48051]= 1284432584;
assign addr[48052]= 1222329801;
assign addr[48053]= 1158676398;
assign addr[48054]= 1093553126;
assign addr[48055]= 1027042599;
assign addr[48056]= 959229189;
assign addr[48057]= 890198924;
assign addr[48058]= 820039373;
assign addr[48059]= 748839539;
assign addr[48060]= 676689746;
assign addr[48061]= 603681519;
assign addr[48062]= 529907477;
assign addr[48063]= 455461206;
assign addr[48064]= 380437148;
assign addr[48065]= 304930476;
assign addr[48066]= 229036977;
assign addr[48067]= 152852926;
assign addr[48068]= 76474970;
assign addr[48069]= 0;
assign addr[48070]= -76474970;
assign addr[48071]= -152852926;
assign addr[48072]= -229036977;
assign addr[48073]= -304930476;
assign addr[48074]= -380437148;
assign addr[48075]= -455461206;
assign addr[48076]= -529907477;
assign addr[48077]= -603681519;
assign addr[48078]= -676689746;
assign addr[48079]= -748839539;
assign addr[48080]= -820039373;
assign addr[48081]= -890198924;
assign addr[48082]= -959229189;
assign addr[48083]= -1027042599;
assign addr[48084]= -1093553126;
assign addr[48085]= -1158676398;
assign addr[48086]= -1222329801;
assign addr[48087]= -1284432584;
assign addr[48088]= -1344905966;
assign addr[48089]= -1403673233;
assign addr[48090]= -1460659832;
assign addr[48091]= -1515793473;
assign addr[48092]= -1569004214;
assign addr[48093]= -1620224553;
assign addr[48094]= -1669389513;
assign addr[48095]= -1716436725;
assign addr[48096]= -1761306505;
assign addr[48097]= -1803941934;
assign addr[48098]= -1844288924;
assign addr[48099]= -1882296293;
assign addr[48100]= -1917915825;
assign addr[48101]= -1951102334;
assign addr[48102]= -1981813720;
assign addr[48103]= -2010011024;
assign addr[48104]= -2035658475;
assign addr[48105]= -2058723538;
assign addr[48106]= -2079176953;
assign addr[48107]= -2096992772;
assign addr[48108]= -2112148396;
assign addr[48109]= -2124624598;
assign addr[48110]= -2134405552;
assign addr[48111]= -2141478848;
assign addr[48112]= -2145835515;
assign addr[48113]= -2147470025;
assign addr[48114]= -2146380306;
assign addr[48115]= -2142567738;
assign addr[48116]= -2136037160;
assign addr[48117]= -2126796855;
assign addr[48118]= -2114858546;
assign addr[48119]= -2100237377;
assign addr[48120]= -2082951896;
assign addr[48121]= -2063024031;
assign addr[48122]= -2040479063;
assign addr[48123]= -2015345591;
assign addr[48124]= -1987655498;
assign addr[48125]= -1957443913;
assign addr[48126]= -1924749160;
assign addr[48127]= -1889612716;
assign addr[48128]= -1852079154;
assign addr[48129]= -1812196087;
assign addr[48130]= -1770014111;
assign addr[48131]= -1725586737;
assign addr[48132]= -1678970324;
assign addr[48133]= -1630224009;
assign addr[48134]= -1579409630;
assign addr[48135]= -1526591649;
assign addr[48136]= -1471837070;
assign addr[48137]= -1415215352;
assign addr[48138]= -1356798326;
assign addr[48139]= -1296660098;
assign addr[48140]= -1234876957;
assign addr[48141]= -1171527280;
assign addr[48142]= -1106691431;
assign addr[48143]= -1040451659;
assign addr[48144]= -972891995;
assign addr[48145]= -904098143;
assign addr[48146]= -834157373;
assign addr[48147]= -763158411;
assign addr[48148]= -691191324;
assign addr[48149]= -618347408;
assign addr[48150]= -544719071;
assign addr[48151]= -470399716;
assign addr[48152]= -395483624;
assign addr[48153]= -320065829;
assign addr[48154]= -244242007;
assign addr[48155]= -168108346;
assign addr[48156]= -91761426;
assign addr[48157]= -15298099;
assign addr[48158]= 61184634;
assign addr[48159]= 137589750;
assign addr[48160]= 213820322;
assign addr[48161]= 289779648;
assign addr[48162]= 365371365;
assign addr[48163]= 440499581;
assign addr[48164]= 515068990;
assign addr[48165]= 588984994;
assign addr[48166]= 662153826;
assign addr[48167]= 734482665;
assign addr[48168]= 805879757;
assign addr[48169]= 876254528;
assign addr[48170]= 945517704;
assign addr[48171]= 1013581418;
assign addr[48172]= 1080359326;
assign addr[48173]= 1145766716;
assign addr[48174]= 1209720613;
assign addr[48175]= 1272139887;
assign addr[48176]= 1332945355;
assign addr[48177]= 1392059879;
assign addr[48178]= 1449408469;
assign addr[48179]= 1504918373;
assign addr[48180]= 1558519173;
assign addr[48181]= 1610142873;
assign addr[48182]= 1659723983;
assign addr[48183]= 1707199606;
assign addr[48184]= 1752509516;
assign addr[48185]= 1795596234;
assign addr[48186]= 1836405100;
assign addr[48187]= 1874884346;
assign addr[48188]= 1910985158;
assign addr[48189]= 1944661739;
assign addr[48190]= 1975871368;
assign addr[48191]= 2004574453;
assign addr[48192]= 2030734582;
assign addr[48193]= 2054318569;
assign addr[48194]= 2075296495;
assign addr[48195]= 2093641749;
assign addr[48196]= 2109331059;
assign addr[48197]= 2122344521;
assign addr[48198]= 2132665626;
assign addr[48199]= 2140281282;
assign addr[48200]= 2145181827;
assign addr[48201]= 2147361045;
assign addr[48202]= 2146816171;
assign addr[48203]= 2143547897;
assign addr[48204]= 2137560369;
assign addr[48205]= 2128861181;
assign addr[48206]= 2117461370;
assign addr[48207]= 2103375398;
assign addr[48208]= 2086621133;
assign addr[48209]= 2067219829;
assign addr[48210]= 2045196100;
assign addr[48211]= 2020577882;
assign addr[48212]= 1993396407;
assign addr[48213]= 1963686155;
assign addr[48214]= 1931484818;
assign addr[48215]= 1896833245;
assign addr[48216]= 1859775393;
assign addr[48217]= 1820358275;
assign addr[48218]= 1778631892;
assign addr[48219]= 1734649179;
assign addr[48220]= 1688465931;
assign addr[48221]= 1640140734;
assign addr[48222]= 1589734894;
assign addr[48223]= 1537312353;
assign addr[48224]= 1482939614;
assign addr[48225]= 1426685652;
assign addr[48226]= 1368621831;
assign addr[48227]= 1308821808;
assign addr[48228]= 1247361445;
assign addr[48229]= 1184318708;
assign addr[48230]= 1119773573;
assign addr[48231]= 1053807919;
assign addr[48232]= 986505429;
assign addr[48233]= 917951481;
assign addr[48234]= 848233042;
assign addr[48235]= 777438554;
assign addr[48236]= 705657826;
assign addr[48237]= 632981917;
assign addr[48238]= 559503022;
assign addr[48239]= 485314355;
assign addr[48240]= 410510029;
assign addr[48241]= 335184940;
assign addr[48242]= 259434643;
assign addr[48243]= 183355234;
assign addr[48244]= 107043224;
assign addr[48245]= 30595422;
assign addr[48246]= -45891193;
assign addr[48247]= -122319591;
assign addr[48248]= -198592817;
assign addr[48249]= -274614114;
assign addr[48250]= -350287041;
assign addr[48251]= -425515602;
assign addr[48252]= -500204365;
assign addr[48253]= -574258580;
assign addr[48254]= -647584304;
assign addr[48255]= -720088517;
assign addr[48256]= -791679244;
assign addr[48257]= -862265664;
assign addr[48258]= -931758235;
assign addr[48259]= -1000068799;
assign addr[48260]= -1067110699;
assign addr[48261]= -1132798888;
assign addr[48262]= -1197050035;
assign addr[48263]= -1259782632;
assign addr[48264]= -1320917099;
assign addr[48265]= -1380375881;
assign addr[48266]= -1438083551;
assign addr[48267]= -1493966902;
assign addr[48268]= -1547955041;
assign addr[48269]= -1599979481;
assign addr[48270]= -1649974225;
assign addr[48271]= -1697875851;
assign addr[48272]= -1743623590;
assign addr[48273]= -1787159411;
assign addr[48274]= -1828428082;
assign addr[48275]= -1867377253;
assign addr[48276]= -1903957513;
assign addr[48277]= -1938122457;
assign addr[48278]= -1969828744;
assign addr[48279]= -1999036154;
assign addr[48280]= -2025707632;
assign addr[48281]= -2049809346;
assign addr[48282]= -2071310720;
assign addr[48283]= -2090184478;
assign addr[48284]= -2106406677;
assign addr[48285]= -2119956737;
assign addr[48286]= -2130817471;
assign addr[48287]= -2138975100;
assign addr[48288]= -2144419275;
assign addr[48289]= -2147143090;
assign addr[48290]= -2147143090;
assign addr[48291]= -2144419275;
assign addr[48292]= -2138975100;
assign addr[48293]= -2130817471;
assign addr[48294]= -2119956737;
assign addr[48295]= -2106406677;
assign addr[48296]= -2090184478;
assign addr[48297]= -2071310720;
assign addr[48298]= -2049809346;
assign addr[48299]= -2025707632;
assign addr[48300]= -1999036154;
assign addr[48301]= -1969828744;
assign addr[48302]= -1938122457;
assign addr[48303]= -1903957513;
assign addr[48304]= -1867377253;
assign addr[48305]= -1828428082;
assign addr[48306]= -1787159411;
assign addr[48307]= -1743623590;
assign addr[48308]= -1697875851;
assign addr[48309]= -1649974225;
assign addr[48310]= -1599979481;
assign addr[48311]= -1547955041;
assign addr[48312]= -1493966902;
assign addr[48313]= -1438083551;
assign addr[48314]= -1380375881;
assign addr[48315]= -1320917099;
assign addr[48316]= -1259782632;
assign addr[48317]= -1197050035;
assign addr[48318]= -1132798888;
assign addr[48319]= -1067110699;
assign addr[48320]= -1000068799;
assign addr[48321]= -931758235;
assign addr[48322]= -862265664;
assign addr[48323]= -791679244;
assign addr[48324]= -720088517;
assign addr[48325]= -647584304;
assign addr[48326]= -574258580;
assign addr[48327]= -500204365;
assign addr[48328]= -425515602;
assign addr[48329]= -350287041;
assign addr[48330]= -274614114;
assign addr[48331]= -198592817;
assign addr[48332]= -122319591;
assign addr[48333]= -45891193;
assign addr[48334]= 30595422;
assign addr[48335]= 107043224;
assign addr[48336]= 183355234;
assign addr[48337]= 259434643;
assign addr[48338]= 335184940;
assign addr[48339]= 410510029;
assign addr[48340]= 485314355;
assign addr[48341]= 559503022;
assign addr[48342]= 632981917;
assign addr[48343]= 705657826;
assign addr[48344]= 777438554;
assign addr[48345]= 848233042;
assign addr[48346]= 917951481;
assign addr[48347]= 986505429;
assign addr[48348]= 1053807919;
assign addr[48349]= 1119773573;
assign addr[48350]= 1184318708;
assign addr[48351]= 1247361445;
assign addr[48352]= 1308821808;
assign addr[48353]= 1368621831;
assign addr[48354]= 1426685652;
assign addr[48355]= 1482939614;
assign addr[48356]= 1537312353;
assign addr[48357]= 1589734894;
assign addr[48358]= 1640140734;
assign addr[48359]= 1688465931;
assign addr[48360]= 1734649179;
assign addr[48361]= 1778631892;
assign addr[48362]= 1820358275;
assign addr[48363]= 1859775393;
assign addr[48364]= 1896833245;
assign addr[48365]= 1931484818;
assign addr[48366]= 1963686155;
assign addr[48367]= 1993396407;
assign addr[48368]= 2020577882;
assign addr[48369]= 2045196100;
assign addr[48370]= 2067219829;
assign addr[48371]= 2086621133;
assign addr[48372]= 2103375398;
assign addr[48373]= 2117461370;
assign addr[48374]= 2128861181;
assign addr[48375]= 2137560369;
assign addr[48376]= 2143547897;
assign addr[48377]= 2146816171;
assign addr[48378]= 2147361045;
assign addr[48379]= 2145181827;
assign addr[48380]= 2140281282;
assign addr[48381]= 2132665626;
assign addr[48382]= 2122344521;
assign addr[48383]= 2109331059;
assign addr[48384]= 2093641749;
assign addr[48385]= 2075296495;
assign addr[48386]= 2054318569;
assign addr[48387]= 2030734582;
assign addr[48388]= 2004574453;
assign addr[48389]= 1975871368;
assign addr[48390]= 1944661739;
assign addr[48391]= 1910985158;
assign addr[48392]= 1874884346;
assign addr[48393]= 1836405100;
assign addr[48394]= 1795596234;
assign addr[48395]= 1752509516;
assign addr[48396]= 1707199606;
assign addr[48397]= 1659723983;
assign addr[48398]= 1610142873;
assign addr[48399]= 1558519173;
assign addr[48400]= 1504918373;
assign addr[48401]= 1449408469;
assign addr[48402]= 1392059879;
assign addr[48403]= 1332945355;
assign addr[48404]= 1272139887;
assign addr[48405]= 1209720613;
assign addr[48406]= 1145766716;
assign addr[48407]= 1080359326;
assign addr[48408]= 1013581418;
assign addr[48409]= 945517704;
assign addr[48410]= 876254528;
assign addr[48411]= 805879757;
assign addr[48412]= 734482665;
assign addr[48413]= 662153826;
assign addr[48414]= 588984994;
assign addr[48415]= 515068990;
assign addr[48416]= 440499581;
assign addr[48417]= 365371365;
assign addr[48418]= 289779648;
assign addr[48419]= 213820322;
assign addr[48420]= 137589750;
assign addr[48421]= 61184634;
assign addr[48422]= -15298099;
assign addr[48423]= -91761426;
assign addr[48424]= -168108346;
assign addr[48425]= -244242007;
assign addr[48426]= -320065829;
assign addr[48427]= -395483624;
assign addr[48428]= -470399716;
assign addr[48429]= -544719071;
assign addr[48430]= -618347408;
assign addr[48431]= -691191324;
assign addr[48432]= -763158411;
assign addr[48433]= -834157373;
assign addr[48434]= -904098143;
assign addr[48435]= -972891995;
assign addr[48436]= -1040451659;
assign addr[48437]= -1106691431;
assign addr[48438]= -1171527280;
assign addr[48439]= -1234876957;
assign addr[48440]= -1296660098;
assign addr[48441]= -1356798326;
assign addr[48442]= -1415215352;
assign addr[48443]= -1471837070;
assign addr[48444]= -1526591649;
assign addr[48445]= -1579409630;
assign addr[48446]= -1630224009;
assign addr[48447]= -1678970324;
assign addr[48448]= -1725586737;
assign addr[48449]= -1770014111;
assign addr[48450]= -1812196087;
assign addr[48451]= -1852079154;
assign addr[48452]= -1889612716;
assign addr[48453]= -1924749160;
assign addr[48454]= -1957443913;
assign addr[48455]= -1987655498;
assign addr[48456]= -2015345591;
assign addr[48457]= -2040479063;
assign addr[48458]= -2063024031;
assign addr[48459]= -2082951896;
assign addr[48460]= -2100237377;
assign addr[48461]= -2114858546;
assign addr[48462]= -2126796855;
assign addr[48463]= -2136037160;
assign addr[48464]= -2142567738;
assign addr[48465]= -2146380306;
assign addr[48466]= -2147470025;
assign addr[48467]= -2145835515;
assign addr[48468]= -2141478848;
assign addr[48469]= -2134405552;
assign addr[48470]= -2124624598;
assign addr[48471]= -2112148396;
assign addr[48472]= -2096992772;
assign addr[48473]= -2079176953;
assign addr[48474]= -2058723538;
assign addr[48475]= -2035658475;
assign addr[48476]= -2010011024;
assign addr[48477]= -1981813720;
assign addr[48478]= -1951102334;
assign addr[48479]= -1917915825;
assign addr[48480]= -1882296293;
assign addr[48481]= -1844288924;
assign addr[48482]= -1803941934;
assign addr[48483]= -1761306505;
assign addr[48484]= -1716436725;
assign addr[48485]= -1669389513;
assign addr[48486]= -1620224553;
assign addr[48487]= -1569004214;
assign addr[48488]= -1515793473;
assign addr[48489]= -1460659832;
assign addr[48490]= -1403673233;
assign addr[48491]= -1344905966;
assign addr[48492]= -1284432584;
assign addr[48493]= -1222329801;
assign addr[48494]= -1158676398;
assign addr[48495]= -1093553126;
assign addr[48496]= -1027042599;
assign addr[48497]= -959229189;
assign addr[48498]= -890198924;
assign addr[48499]= -820039373;
assign addr[48500]= -748839539;
assign addr[48501]= -676689746;
assign addr[48502]= -603681519;
assign addr[48503]= -529907477;
assign addr[48504]= -455461206;
assign addr[48505]= -380437148;
assign addr[48506]= -304930476;
assign addr[48507]= -229036977;
assign addr[48508]= -152852926;
assign addr[48509]= -76474970;
assign addr[48510]= 0;
assign addr[48511]= 76474970;
assign addr[48512]= 152852926;
assign addr[48513]= 229036977;
assign addr[48514]= 304930476;
assign addr[48515]= 380437148;
assign addr[48516]= 455461206;
assign addr[48517]= 529907477;
assign addr[48518]= 603681519;
assign addr[48519]= 676689746;
assign addr[48520]= 748839539;
assign addr[48521]= 820039373;
assign addr[48522]= 890198924;
assign addr[48523]= 959229189;
assign addr[48524]= 1027042599;
assign addr[48525]= 1093553126;
assign addr[48526]= 1158676398;
assign addr[48527]= 1222329801;
assign addr[48528]= 1284432584;
assign addr[48529]= 1344905966;
assign addr[48530]= 1403673233;
assign addr[48531]= 1460659832;
assign addr[48532]= 1515793473;
assign addr[48533]= 1569004214;
assign addr[48534]= 1620224553;
assign addr[48535]= 1669389513;
assign addr[48536]= 1716436725;
assign addr[48537]= 1761306505;
assign addr[48538]= 1803941934;
assign addr[48539]= 1844288924;
assign addr[48540]= 1882296293;
assign addr[48541]= 1917915825;
assign addr[48542]= 1951102334;
assign addr[48543]= 1981813720;
assign addr[48544]= 2010011024;
assign addr[48545]= 2035658475;
assign addr[48546]= 2058723538;
assign addr[48547]= 2079176953;
assign addr[48548]= 2096992772;
assign addr[48549]= 2112148396;
assign addr[48550]= 2124624598;
assign addr[48551]= 2134405552;
assign addr[48552]= 2141478848;
assign addr[48553]= 2145835515;
assign addr[48554]= 2147470025;
assign addr[48555]= 2146380306;
assign addr[48556]= 2142567738;
assign addr[48557]= 2136037160;
assign addr[48558]= 2126796855;
assign addr[48559]= 2114858546;
assign addr[48560]= 2100237377;
assign addr[48561]= 2082951896;
assign addr[48562]= 2063024031;
assign addr[48563]= 2040479063;
assign addr[48564]= 2015345591;
assign addr[48565]= 1987655498;
assign addr[48566]= 1957443913;
assign addr[48567]= 1924749160;
assign addr[48568]= 1889612716;
assign addr[48569]= 1852079154;
assign addr[48570]= 1812196087;
assign addr[48571]= 1770014111;
assign addr[48572]= 1725586737;
assign addr[48573]= 1678970324;
assign addr[48574]= 1630224009;
assign addr[48575]= 1579409630;
assign addr[48576]= 1526591649;
assign addr[48577]= 1471837070;
assign addr[48578]= 1415215352;
assign addr[48579]= 1356798326;
assign addr[48580]= 1296660098;
assign addr[48581]= 1234876957;
assign addr[48582]= 1171527280;
assign addr[48583]= 1106691431;
assign addr[48584]= 1040451659;
assign addr[48585]= 972891995;
assign addr[48586]= 904098143;
assign addr[48587]= 834157373;
assign addr[48588]= 763158411;
assign addr[48589]= 691191324;
assign addr[48590]= 618347408;
assign addr[48591]= 544719071;
assign addr[48592]= 470399716;
assign addr[48593]= 395483624;
assign addr[48594]= 320065829;
assign addr[48595]= 244242007;
assign addr[48596]= 168108346;
assign addr[48597]= 91761426;
assign addr[48598]= 15298099;
assign addr[48599]= -61184634;
assign addr[48600]= -137589750;
assign addr[48601]= -213820322;
assign addr[48602]= -289779648;
assign addr[48603]= -365371365;
assign addr[48604]= -440499581;
assign addr[48605]= -515068990;
assign addr[48606]= -588984994;
assign addr[48607]= -662153826;
assign addr[48608]= -734482665;
assign addr[48609]= -805879757;
assign addr[48610]= -876254528;
assign addr[48611]= -945517704;
assign addr[48612]= -1013581418;
assign addr[48613]= -1080359326;
assign addr[48614]= -1145766716;
assign addr[48615]= -1209720613;
assign addr[48616]= -1272139887;
assign addr[48617]= -1332945355;
assign addr[48618]= -1392059879;
assign addr[48619]= -1449408469;
assign addr[48620]= -1504918373;
assign addr[48621]= -1558519173;
assign addr[48622]= -1610142873;
assign addr[48623]= -1659723983;
assign addr[48624]= -1707199606;
assign addr[48625]= -1752509516;
assign addr[48626]= -1795596234;
assign addr[48627]= -1836405100;
assign addr[48628]= -1874884346;
assign addr[48629]= -1910985158;
assign addr[48630]= -1944661739;
assign addr[48631]= -1975871368;
assign addr[48632]= -2004574453;
assign addr[48633]= -2030734582;
assign addr[48634]= -2054318569;
assign addr[48635]= -2075296495;
assign addr[48636]= -2093641749;
assign addr[48637]= -2109331059;
assign addr[48638]= -2122344521;
assign addr[48639]= -2132665626;
assign addr[48640]= -2140281282;
assign addr[48641]= -2145181827;
assign addr[48642]= -2147361045;
assign addr[48643]= -2146816171;
assign addr[48644]= -2143547897;
assign addr[48645]= -2137560369;
assign addr[48646]= -2128861181;
assign addr[48647]= -2117461370;
assign addr[48648]= -2103375398;
assign addr[48649]= -2086621133;
assign addr[48650]= -2067219829;
assign addr[48651]= -2045196100;
assign addr[48652]= -2020577882;
assign addr[48653]= -1993396407;
assign addr[48654]= -1963686155;
assign addr[48655]= -1931484818;
assign addr[48656]= -1896833245;
assign addr[48657]= -1859775393;
assign addr[48658]= -1820358275;
assign addr[48659]= -1778631892;
assign addr[48660]= -1734649179;
assign addr[48661]= -1688465931;
assign addr[48662]= -1640140734;
assign addr[48663]= -1589734894;
assign addr[48664]= -1537312353;
assign addr[48665]= -1482939614;
assign addr[48666]= -1426685652;
assign addr[48667]= -1368621831;
assign addr[48668]= -1308821808;
assign addr[48669]= -1247361445;
assign addr[48670]= -1184318708;
assign addr[48671]= -1119773573;
assign addr[48672]= -1053807919;
assign addr[48673]= -986505429;
assign addr[48674]= -917951481;
assign addr[48675]= -848233042;
assign addr[48676]= -777438554;
assign addr[48677]= -705657826;
assign addr[48678]= -632981917;
assign addr[48679]= -559503022;
assign addr[48680]= -485314355;
assign addr[48681]= -410510029;
assign addr[48682]= -335184940;
assign addr[48683]= -259434643;
assign addr[48684]= -183355234;
assign addr[48685]= -107043224;
assign addr[48686]= -30595422;
assign addr[48687]= 45891193;
assign addr[48688]= 122319591;
assign addr[48689]= 198592817;
assign addr[48690]= 274614114;
assign addr[48691]= 350287041;
assign addr[48692]= 425515602;
assign addr[48693]= 500204365;
assign addr[48694]= 574258580;
assign addr[48695]= 647584304;
assign addr[48696]= 720088517;
assign addr[48697]= 791679244;
assign addr[48698]= 862265664;
assign addr[48699]= 931758235;
assign addr[48700]= 1000068799;
assign addr[48701]= 1067110699;
assign addr[48702]= 1132798888;
assign addr[48703]= 1197050035;
assign addr[48704]= 1259782632;
assign addr[48705]= 1320917099;
assign addr[48706]= 1380375881;
assign addr[48707]= 1438083551;
assign addr[48708]= 1493966902;
assign addr[48709]= 1547955041;
assign addr[48710]= 1599979481;
assign addr[48711]= 1649974225;
assign addr[48712]= 1697875851;
assign addr[48713]= 1743623590;
assign addr[48714]= 1787159411;
assign addr[48715]= 1828428082;
assign addr[48716]= 1867377253;
assign addr[48717]= 1903957513;
assign addr[48718]= 1938122457;
assign addr[48719]= 1969828744;
assign addr[48720]= 1999036154;
assign addr[48721]= 2025707632;
assign addr[48722]= 2049809346;
assign addr[48723]= 2071310720;
assign addr[48724]= 2090184478;
assign addr[48725]= 2106406677;
assign addr[48726]= 2119956737;
assign addr[48727]= 2130817471;
assign addr[48728]= 2138975100;
assign addr[48729]= 2144419275;
assign addr[48730]= 2147143090;
assign addr[48731]= 2147143090;
assign addr[48732]= 2144419275;
assign addr[48733]= 2138975100;
assign addr[48734]= 2130817471;
assign addr[48735]= 2119956737;
assign addr[48736]= 2106406677;
assign addr[48737]= 2090184478;
assign addr[48738]= 2071310720;
assign addr[48739]= 2049809346;
assign addr[48740]= 2025707632;
assign addr[48741]= 1999036154;
assign addr[48742]= 1969828744;
assign addr[48743]= 1938122457;
assign addr[48744]= 1903957513;
assign addr[48745]= 1867377253;
assign addr[48746]= 1828428082;
assign addr[48747]= 1787159411;
assign addr[48748]= 1743623590;
assign addr[48749]= 1697875851;
assign addr[48750]= 1649974225;
assign addr[48751]= 1599979481;
assign addr[48752]= 1547955041;
assign addr[48753]= 1493966902;
assign addr[48754]= 1438083551;
assign addr[48755]= 1380375881;
assign addr[48756]= 1320917099;
assign addr[48757]= 1259782632;
assign addr[48758]= 1197050035;
assign addr[48759]= 1132798888;
assign addr[48760]= 1067110699;
assign addr[48761]= 1000068799;
assign addr[48762]= 931758235;
assign addr[48763]= 862265664;
assign addr[48764]= 791679244;
assign addr[48765]= 720088517;
assign addr[48766]= 647584304;
assign addr[48767]= 574258580;
assign addr[48768]= 500204365;
assign addr[48769]= 425515602;
assign addr[48770]= 350287041;
assign addr[48771]= 274614114;
assign addr[48772]= 198592817;
assign addr[48773]= 122319591;
assign addr[48774]= 45891193;
assign addr[48775]= -30595422;
assign addr[48776]= -107043224;
assign addr[48777]= -183355234;
assign addr[48778]= -259434643;
assign addr[48779]= -335184940;
assign addr[48780]= -410510029;
assign addr[48781]= -485314355;
assign addr[48782]= -559503022;
assign addr[48783]= -632981917;
assign addr[48784]= -705657826;
assign addr[48785]= -777438554;
assign addr[48786]= -848233042;
assign addr[48787]= -917951481;
assign addr[48788]= -986505429;
assign addr[48789]= -1053807919;
assign addr[48790]= -1119773573;
assign addr[48791]= -1184318708;
assign addr[48792]= -1247361445;
assign addr[48793]= -1308821808;
assign addr[48794]= -1368621831;
assign addr[48795]= -1426685652;
assign addr[48796]= -1482939614;
assign addr[48797]= -1537312353;
assign addr[48798]= -1589734894;
assign addr[48799]= -1640140734;
assign addr[48800]= -1688465931;
assign addr[48801]= -1734649179;
assign addr[48802]= -1778631892;
assign addr[48803]= -1820358275;
assign addr[48804]= -1859775393;
assign addr[48805]= -1896833245;
assign addr[48806]= -1931484818;
assign addr[48807]= -1963686155;
assign addr[48808]= -1993396407;
assign addr[48809]= -2020577882;
assign addr[48810]= -2045196100;
assign addr[48811]= -2067219829;
assign addr[48812]= -2086621133;
assign addr[48813]= -2103375398;
assign addr[48814]= -2117461370;
assign addr[48815]= -2128861181;
assign addr[48816]= -2137560369;
assign addr[48817]= -2143547897;
assign addr[48818]= -2146816171;
assign addr[48819]= -2147361045;
assign addr[48820]= -2145181827;
assign addr[48821]= -2140281282;
assign addr[48822]= -2132665626;
assign addr[48823]= -2122344521;
assign addr[48824]= -2109331059;
assign addr[48825]= -2093641749;
assign addr[48826]= -2075296495;
assign addr[48827]= -2054318569;
assign addr[48828]= -2030734582;
assign addr[48829]= -2004574453;
assign addr[48830]= -1975871368;
assign addr[48831]= -1944661739;
assign addr[48832]= -1910985158;
assign addr[48833]= -1874884346;
assign addr[48834]= -1836405100;
assign addr[48835]= -1795596234;
assign addr[48836]= -1752509516;
assign addr[48837]= -1707199606;
assign addr[48838]= -1659723983;
assign addr[48839]= -1610142873;
assign addr[48840]= -1558519173;
assign addr[48841]= -1504918373;
assign addr[48842]= -1449408469;
assign addr[48843]= -1392059879;
assign addr[48844]= -1332945355;
assign addr[48845]= -1272139887;
assign addr[48846]= -1209720613;
assign addr[48847]= -1145766716;
assign addr[48848]= -1080359326;
assign addr[48849]= -1013581418;
assign addr[48850]= -945517704;
assign addr[48851]= -876254528;
assign addr[48852]= -805879757;
assign addr[48853]= -734482665;
assign addr[48854]= -662153826;
assign addr[48855]= -588984994;
assign addr[48856]= -515068990;
assign addr[48857]= -440499581;
assign addr[48858]= -365371365;
assign addr[48859]= -289779648;
assign addr[48860]= -213820322;
assign addr[48861]= -137589750;
assign addr[48862]= -61184634;
assign addr[48863]= 15298099;
assign addr[48864]= 91761426;
assign addr[48865]= 168108346;
assign addr[48866]= 244242007;
assign addr[48867]= 320065829;
assign addr[48868]= 395483624;
assign addr[48869]= 470399716;
assign addr[48870]= 544719071;
assign addr[48871]= 618347408;
assign addr[48872]= 691191324;
assign addr[48873]= 763158411;
assign addr[48874]= 834157373;
assign addr[48875]= 904098143;
assign addr[48876]= 972891995;
assign addr[48877]= 1040451659;
assign addr[48878]= 1106691431;
assign addr[48879]= 1171527280;
assign addr[48880]= 1234876957;
assign addr[48881]= 1296660098;
assign addr[48882]= 1356798326;
assign addr[48883]= 1415215352;
assign addr[48884]= 1471837070;
assign addr[48885]= 1526591649;
assign addr[48886]= 1579409630;
assign addr[48887]= 1630224009;
assign addr[48888]= 1678970324;
assign addr[48889]= 1725586737;
assign addr[48890]= 1770014111;
assign addr[48891]= 1812196087;
assign addr[48892]= 1852079154;
assign addr[48893]= 1889612716;
assign addr[48894]= 1924749160;
assign addr[48895]= 1957443913;
assign addr[48896]= 1987655498;
assign addr[48897]= 2015345591;
assign addr[48898]= 2040479063;
assign addr[48899]= 2063024031;
assign addr[48900]= 2082951896;
assign addr[48901]= 2100237377;
assign addr[48902]= 2114858546;
assign addr[48903]= 2126796855;
assign addr[48904]= 2136037160;
assign addr[48905]= 2142567738;
assign addr[48906]= 2146380306;
assign addr[48907]= 2147470025;
assign addr[48908]= 2145835515;
assign addr[48909]= 2141478848;
assign addr[48910]= 2134405552;
assign addr[48911]= 2124624598;
assign addr[48912]= 2112148396;
assign addr[48913]= 2096992772;
assign addr[48914]= 2079176953;
assign addr[48915]= 2058723538;
assign addr[48916]= 2035658475;
assign addr[48917]= 2010011024;
assign addr[48918]= 1981813720;
assign addr[48919]= 1951102334;
assign addr[48920]= 1917915825;
assign addr[48921]= 1882296293;
assign addr[48922]= 1844288924;
assign addr[48923]= 1803941934;
assign addr[48924]= 1761306505;
assign addr[48925]= 1716436725;
assign addr[48926]= 1669389513;
assign addr[48927]= 1620224553;
assign addr[48928]= 1569004214;
assign addr[48929]= 1515793473;
assign addr[48930]= 1460659832;
assign addr[48931]= 1403673233;
assign addr[48932]= 1344905966;
assign addr[48933]= 1284432584;
assign addr[48934]= 1222329801;
assign addr[48935]= 1158676398;
assign addr[48936]= 1093553126;
assign addr[48937]= 1027042599;
assign addr[48938]= 959229189;
assign addr[48939]= 890198924;
assign addr[48940]= 820039373;
assign addr[48941]= 748839539;
assign addr[48942]= 676689746;
assign addr[48943]= 603681519;
assign addr[48944]= 529907477;
assign addr[48945]= 455461206;
assign addr[48946]= 380437148;
assign addr[48947]= 304930476;
assign addr[48948]= 229036977;
assign addr[48949]= 152852926;
assign addr[48950]= 76474970;
assign addr[48951]= 0;
assign addr[48952]= -76474970;
assign addr[48953]= -152852926;
assign addr[48954]= -229036977;
assign addr[48955]= -304930476;
assign addr[48956]= -380437148;
assign addr[48957]= -455461206;
assign addr[48958]= -529907477;
assign addr[48959]= -603681519;
assign addr[48960]= -676689746;
assign addr[48961]= -748839539;
assign addr[48962]= -820039373;
assign addr[48963]= -890198924;
assign addr[48964]= -959229189;
assign addr[48965]= -1027042599;
assign addr[48966]= -1093553126;
assign addr[48967]= -1158676398;
assign addr[48968]= -1222329801;
assign addr[48969]= -1284432584;
assign addr[48970]= -1344905966;
assign addr[48971]= -1403673233;
assign addr[48972]= -1460659832;
assign addr[48973]= -1515793473;
assign addr[48974]= -1569004214;
assign addr[48975]= -1620224553;
assign addr[48976]= -1669389513;
assign addr[48977]= -1716436725;
assign addr[48978]= -1761306505;
assign addr[48979]= -1803941934;
assign addr[48980]= -1844288924;
assign addr[48981]= -1882296293;
assign addr[48982]= -1917915825;
assign addr[48983]= -1951102334;
assign addr[48984]= -1981813720;
assign addr[48985]= -2010011024;
assign addr[48986]= -2035658475;
assign addr[48987]= -2058723538;
assign addr[48988]= -2079176953;
assign addr[48989]= -2096992772;
assign addr[48990]= -2112148396;
assign addr[48991]= -2124624598;
assign addr[48992]= -2134405552;
assign addr[48993]= -2141478848;
assign addr[48994]= -2145835515;
assign addr[48995]= -2147470025;
assign addr[48996]= -2146380306;
assign addr[48997]= -2142567738;
assign addr[48998]= -2136037160;
assign addr[48999]= -2126796855;
assign addr[49000]= -2114858546;
assign addr[49001]= -2100237377;
assign addr[49002]= -2082951896;
assign addr[49003]= -2063024031;
assign addr[49004]= -2040479063;
assign addr[49005]= -2015345591;
assign addr[49006]= -1987655498;
assign addr[49007]= -1957443913;
assign addr[49008]= -1924749160;
assign addr[49009]= -1889612716;
assign addr[49010]= -1852079154;
assign addr[49011]= -1812196087;
assign addr[49012]= -1770014111;
assign addr[49013]= -1725586737;
assign addr[49014]= -1678970324;
assign addr[49015]= -1630224009;
assign addr[49016]= -1579409630;
assign addr[49017]= -1526591649;
assign addr[49018]= -1471837070;
assign addr[49019]= -1415215352;
assign addr[49020]= -1356798326;
assign addr[49021]= -1296660098;
assign addr[49022]= -1234876957;
assign addr[49023]= -1171527280;
assign addr[49024]= -1106691431;
assign addr[49025]= -1040451659;
assign addr[49026]= -972891995;
assign addr[49027]= -904098143;
assign addr[49028]= -834157373;
assign addr[49029]= -763158411;
assign addr[49030]= -691191324;
assign addr[49031]= -618347408;
assign addr[49032]= -544719071;
assign addr[49033]= -470399716;
assign addr[49034]= -395483624;
assign addr[49035]= -320065829;
assign addr[49036]= -244242007;
assign addr[49037]= -168108346;
assign addr[49038]= -91761426;
assign addr[49039]= -15298099;
assign addr[49040]= 61184634;
assign addr[49041]= 137589750;
assign addr[49042]= 213820322;
assign addr[49043]= 289779648;
assign addr[49044]= 365371365;
assign addr[49045]= 440499581;
assign addr[49046]= 515068990;
assign addr[49047]= 588984994;
assign addr[49048]= 662153826;
assign addr[49049]= 734482665;
assign addr[49050]= 805879757;
assign addr[49051]= 876254528;
assign addr[49052]= 945517704;
assign addr[49053]= 1013581418;
assign addr[49054]= 1080359326;
assign addr[49055]= 1145766716;
assign addr[49056]= 1209720613;
assign addr[49057]= 1272139887;
assign addr[49058]= 1332945355;
assign addr[49059]= 1392059879;
assign addr[49060]= 1449408469;
assign addr[49061]= 1504918373;
assign addr[49062]= 1558519173;
assign addr[49063]= 1610142873;
assign addr[49064]= 1659723983;
assign addr[49065]= 1707199606;
assign addr[49066]= 1752509516;
assign addr[49067]= 1795596234;
assign addr[49068]= 1836405100;
assign addr[49069]= 1874884346;
assign addr[49070]= 1910985158;
assign addr[49071]= 1944661739;
assign addr[49072]= 1975871368;
assign addr[49073]= 2004574453;
assign addr[49074]= 2030734582;
assign addr[49075]= 2054318569;
assign addr[49076]= 2075296495;
assign addr[49077]= 2093641749;
assign addr[49078]= 2109331059;
assign addr[49079]= 2122344521;
assign addr[49080]= 2132665626;
assign addr[49081]= 2140281282;
assign addr[49082]= 2145181827;
assign addr[49083]= 2147361045;
assign addr[49084]= 2146816171;
assign addr[49085]= 2143547897;
assign addr[49086]= 2137560369;
assign addr[49087]= 2128861181;
assign addr[49088]= 2117461370;
assign addr[49089]= 2103375398;
assign addr[49090]= 2086621133;
assign addr[49091]= 2067219829;
assign addr[49092]= 2045196100;
assign addr[49093]= 2020577882;
assign addr[49094]= 1993396407;
assign addr[49095]= 1963686155;
assign addr[49096]= 1931484818;
assign addr[49097]= 1896833245;
assign addr[49098]= 1859775393;
assign addr[49099]= 1820358275;
assign addr[49100]= 1778631892;
assign addr[49101]= 1734649179;
assign addr[49102]= 1688465931;
assign addr[49103]= 1640140734;
assign addr[49104]= 1589734894;
assign addr[49105]= 1537312353;
assign addr[49106]= 1482939614;
assign addr[49107]= 1426685652;
assign addr[49108]= 1368621831;
assign addr[49109]= 1308821808;
assign addr[49110]= 1247361445;
assign addr[49111]= 1184318708;
assign addr[49112]= 1119773573;
assign addr[49113]= 1053807919;
assign addr[49114]= 986505429;
assign addr[49115]= 917951481;
assign addr[49116]= 848233042;
assign addr[49117]= 777438554;
assign addr[49118]= 705657826;
assign addr[49119]= 632981917;
assign addr[49120]= 559503022;
assign addr[49121]= 485314355;
assign addr[49122]= 410510029;
assign addr[49123]= 335184940;
assign addr[49124]= 259434643;
assign addr[49125]= 183355234;
assign addr[49126]= 107043224;
assign addr[49127]= 30595422;
assign addr[49128]= -45891193;
assign addr[49129]= -122319591;
assign addr[49130]= -198592817;
assign addr[49131]= -274614114;
assign addr[49132]= -350287041;
assign addr[49133]= -425515602;
assign addr[49134]= -500204365;
assign addr[49135]= -574258580;
assign addr[49136]= -647584304;
assign addr[49137]= -720088517;
assign addr[49138]= -791679244;
assign addr[49139]= -862265664;
assign addr[49140]= -931758235;
assign addr[49141]= -1000068799;
assign addr[49142]= -1067110699;
assign addr[49143]= -1132798888;
assign addr[49144]= -1197050035;
assign addr[49145]= -1259782632;
assign addr[49146]= -1320917099;
assign addr[49147]= -1380375881;
assign addr[49148]= -1438083551;
assign addr[49149]= -1493966902;
assign addr[49150]= -1547955041;
assign addr[49151]= -1599979481;
assign addr[49152]= -1649974225;
assign addr[49153]= -1697875851;
assign addr[49154]= -1743623590;
assign addr[49155]= -1787159411;
assign addr[49156]= -1828428082;
assign addr[49157]= -1867377253;
assign addr[49158]= -1903957513;
assign addr[49159]= -1938122457;
assign addr[49160]= -1969828744;
assign addr[49161]= -1999036154;
assign addr[49162]= -2025707632;
assign addr[49163]= -2049809346;
assign addr[49164]= -2071310720;
assign addr[49165]= -2090184478;
assign addr[49166]= -2106406677;
assign addr[49167]= -2119956737;
assign addr[49168]= -2130817471;
assign addr[49169]= -2138975100;
assign addr[49170]= -2144419275;
assign addr[49171]= -2147143090;
assign addr[49172]= -2147143090;
assign addr[49173]= -2144419275;
assign addr[49174]= -2138975100;
assign addr[49175]= -2130817471;
assign addr[49176]= -2119956737;
assign addr[49177]= -2106406677;
assign addr[49178]= -2090184478;
assign addr[49179]= -2071310720;
assign addr[49180]= -2049809346;
assign addr[49181]= -2025707632;
assign addr[49182]= -1999036154;
assign addr[49183]= -1969828744;
assign addr[49184]= -1938122457;
assign addr[49185]= -1903957513;
assign addr[49186]= -1867377253;
assign addr[49187]= -1828428082;
assign addr[49188]= -1787159411;
assign addr[49189]= -1743623590;
assign addr[49190]= -1697875851;
assign addr[49191]= -1649974225;
assign addr[49192]= -1599979481;
assign addr[49193]= -1547955041;
assign addr[49194]= -1493966902;
assign addr[49195]= -1438083551;
assign addr[49196]= -1380375881;
assign addr[49197]= -1320917099;
assign addr[49198]= -1259782632;
assign addr[49199]= -1197050035;
assign addr[49200]= -1132798888;
assign addr[49201]= -1067110699;
assign addr[49202]= -1000068799;
assign addr[49203]= -931758235;
assign addr[49204]= -862265664;
assign addr[49205]= -791679244;
assign addr[49206]= -720088517;
assign addr[49207]= -647584304;
assign addr[49208]= -574258580;
assign addr[49209]= -500204365;
assign addr[49210]= -425515602;
assign addr[49211]= -350287041;
assign addr[49212]= -274614114;
assign addr[49213]= -198592817;
assign addr[49214]= -122319591;
assign addr[49215]= -45891193;
assign addr[49216]= 30595422;
assign addr[49217]= 107043224;
assign addr[49218]= 183355234;
assign addr[49219]= 259434643;
assign addr[49220]= 335184940;
assign addr[49221]= 410510029;
assign addr[49222]= 485314355;
assign addr[49223]= 559503022;
assign addr[49224]= 632981917;
assign addr[49225]= 705657826;
assign addr[49226]= 777438554;
assign addr[49227]= 848233042;
assign addr[49228]= 917951481;
assign addr[49229]= 986505429;
assign addr[49230]= 1053807919;
assign addr[49231]= 1119773573;
assign addr[49232]= 1184318708;
assign addr[49233]= 1247361445;
assign addr[49234]= 1308821808;
assign addr[49235]= 1368621831;
assign addr[49236]= 1426685652;
assign addr[49237]= 1482939614;
assign addr[49238]= 1537312353;
assign addr[49239]= 1589734894;
assign addr[49240]= 1640140734;
assign addr[49241]= 1688465931;
assign addr[49242]= 1734649179;
assign addr[49243]= 1778631892;
assign addr[49244]= 1820358275;
assign addr[49245]= 1859775393;
assign addr[49246]= 1896833245;
assign addr[49247]= 1931484818;
assign addr[49248]= 1963686155;
assign addr[49249]= 1993396407;
assign addr[49250]= 2020577882;
assign addr[49251]= 2045196100;
assign addr[49252]= 2067219829;
assign addr[49253]= 2086621133;
assign addr[49254]= 2103375398;
assign addr[49255]= 2117461370;
assign addr[49256]= 2128861181;
assign addr[49257]= 2137560369;
assign addr[49258]= 2143547897;
assign addr[49259]= 2146816171;
assign addr[49260]= 2147361045;
assign addr[49261]= 2145181827;
assign addr[49262]= 2140281282;
assign addr[49263]= 2132665626;
assign addr[49264]= 2122344521;
assign addr[49265]= 2109331059;
assign addr[49266]= 2093641749;
assign addr[49267]= 2075296495;
assign addr[49268]= 2054318569;
assign addr[49269]= 2030734582;
assign addr[49270]= 2004574453;
assign addr[49271]= 1975871368;
assign addr[49272]= 1944661739;
assign addr[49273]= 1910985158;
assign addr[49274]= 1874884346;
assign addr[49275]= 1836405100;
assign addr[49276]= 1795596234;
assign addr[49277]= 1752509516;
assign addr[49278]= 1707199606;
assign addr[49279]= 1659723983;
assign addr[49280]= 1610142873;
assign addr[49281]= 1558519173;
assign addr[49282]= 1504918373;
assign addr[49283]= 1449408469;
assign addr[49284]= 1392059879;
assign addr[49285]= 1332945355;
assign addr[49286]= 1272139887;
assign addr[49287]= 1209720613;
assign addr[49288]= 1145766716;
assign addr[49289]= 1080359326;
assign addr[49290]= 1013581418;
assign addr[49291]= 945517704;
assign addr[49292]= 876254528;
assign addr[49293]= 805879757;
assign addr[49294]= 734482665;
assign addr[49295]= 662153826;
assign addr[49296]= 588984994;
assign addr[49297]= 515068990;
assign addr[49298]= 440499581;
assign addr[49299]= 365371365;
assign addr[49300]= 289779648;
assign addr[49301]= 213820322;
assign addr[49302]= 137589750;
assign addr[49303]= 61184634;
assign addr[49304]= -15298099;
assign addr[49305]= -91761426;
assign addr[49306]= -168108346;
assign addr[49307]= -244242007;
assign addr[49308]= -320065829;
assign addr[49309]= -395483624;
assign addr[49310]= -470399716;
assign addr[49311]= -544719071;
assign addr[49312]= -618347408;
assign addr[49313]= -691191324;
assign addr[49314]= -763158411;
assign addr[49315]= -834157373;
assign addr[49316]= -904098143;
assign addr[49317]= -972891995;
assign addr[49318]= -1040451659;
assign addr[49319]= -1106691431;
assign addr[49320]= -1171527280;
assign addr[49321]= -1234876957;
assign addr[49322]= -1296660098;
assign addr[49323]= -1356798326;
assign addr[49324]= -1415215352;
assign addr[49325]= -1471837070;
assign addr[49326]= -1526591649;
assign addr[49327]= -1579409630;
assign addr[49328]= -1630224009;
assign addr[49329]= -1678970324;
assign addr[49330]= -1725586737;
assign addr[49331]= -1770014111;
assign addr[49332]= -1812196087;
assign addr[49333]= -1852079154;
assign addr[49334]= -1889612716;
assign addr[49335]= -1924749160;
assign addr[49336]= -1957443913;
assign addr[49337]= -1987655498;
assign addr[49338]= -2015345591;
assign addr[49339]= -2040479063;
assign addr[49340]= -2063024031;
assign addr[49341]= -2082951896;
assign addr[49342]= -2100237377;
assign addr[49343]= -2114858546;
assign addr[49344]= -2126796855;
assign addr[49345]= -2136037160;
assign addr[49346]= -2142567738;
assign addr[49347]= -2146380306;
assign addr[49348]= -2147470025;
assign addr[49349]= -2145835515;
assign addr[49350]= -2141478848;
assign addr[49351]= -2134405552;
assign addr[49352]= -2124624598;
assign addr[49353]= -2112148396;
assign addr[49354]= -2096992772;
assign addr[49355]= -2079176953;
assign addr[49356]= -2058723538;
assign addr[49357]= -2035658475;
assign addr[49358]= -2010011024;
assign addr[49359]= -1981813720;
assign addr[49360]= -1951102334;
assign addr[49361]= -1917915825;
assign addr[49362]= -1882296293;
assign addr[49363]= -1844288924;
assign addr[49364]= -1803941934;
assign addr[49365]= -1761306505;
assign addr[49366]= -1716436725;
assign addr[49367]= -1669389513;
assign addr[49368]= -1620224553;
assign addr[49369]= -1569004214;
assign addr[49370]= -1515793473;
assign addr[49371]= -1460659832;
assign addr[49372]= -1403673233;
assign addr[49373]= -1344905966;
assign addr[49374]= -1284432584;
assign addr[49375]= -1222329801;
assign addr[49376]= -1158676398;
assign addr[49377]= -1093553126;
assign addr[49378]= -1027042599;
assign addr[49379]= -959229189;
assign addr[49380]= -890198924;
assign addr[49381]= -820039373;
assign addr[49382]= -748839539;
assign addr[49383]= -676689746;
assign addr[49384]= -603681519;
assign addr[49385]= -529907477;
assign addr[49386]= -455461206;
assign addr[49387]= -380437148;
assign addr[49388]= -304930476;
assign addr[49389]= -229036977;
assign addr[49390]= -152852926;
assign addr[49391]= -76474970;
assign addr[49392]= 0;
assign addr[49393]= 76474970;
assign addr[49394]= 152852926;
assign addr[49395]= 229036977;
assign addr[49396]= 304930476;
assign addr[49397]= 380437148;
assign addr[49398]= 455461206;
assign addr[49399]= 529907477;
assign addr[49400]= 603681519;
assign addr[49401]= 676689746;
assign addr[49402]= 748839539;
assign addr[49403]= 820039373;
assign addr[49404]= 890198924;
assign addr[49405]= 959229189;
assign addr[49406]= 1027042599;
assign addr[49407]= 1093553126;
assign addr[49408]= 1158676398;
assign addr[49409]= 1222329801;
assign addr[49410]= 1284432584;
assign addr[49411]= 1344905966;
assign addr[49412]= 1403673233;
assign addr[49413]= 1460659832;
assign addr[49414]= 1515793473;
assign addr[49415]= 1569004214;
assign addr[49416]= 1620224553;
assign addr[49417]= 1669389513;
assign addr[49418]= 1716436725;
assign addr[49419]= 1761306505;
assign addr[49420]= 1803941934;
assign addr[49421]= 1844288924;
assign addr[49422]= 1882296293;
assign addr[49423]= 1917915825;
assign addr[49424]= 1951102334;
assign addr[49425]= 1981813720;
assign addr[49426]= 2010011024;
assign addr[49427]= 2035658475;
assign addr[49428]= 2058723538;
assign addr[49429]= 2079176953;
assign addr[49430]= 2096992772;
assign addr[49431]= 2112148396;
assign addr[49432]= 2124624598;
assign addr[49433]= 2134405552;
assign addr[49434]= 2141478848;
assign addr[49435]= 2145835515;
assign addr[49436]= 2147470025;
assign addr[49437]= 2146380306;
assign addr[49438]= 2142567738;
assign addr[49439]= 2136037160;
assign addr[49440]= 2126796855;
assign addr[49441]= 2114858546;
assign addr[49442]= 2100237377;
assign addr[49443]= 2082951896;
assign addr[49444]= 2063024031;
assign addr[49445]= 2040479063;
assign addr[49446]= 2015345591;
assign addr[49447]= 1987655498;
assign addr[49448]= 1957443913;
assign addr[49449]= 1924749160;
assign addr[49450]= 1889612716;
assign addr[49451]= 1852079154;
assign addr[49452]= 1812196087;
assign addr[49453]= 1770014111;
assign addr[49454]= 1725586737;
assign addr[49455]= 1678970324;
assign addr[49456]= 1630224009;
assign addr[49457]= 1579409630;
assign addr[49458]= 1526591649;
assign addr[49459]= 1471837070;
assign addr[49460]= 1415215352;
assign addr[49461]= 1356798326;
assign addr[49462]= 1296660098;
assign addr[49463]= 1234876957;
assign addr[49464]= 1171527280;
assign addr[49465]= 1106691431;
assign addr[49466]= 1040451659;
assign addr[49467]= 972891995;
assign addr[49468]= 904098143;
assign addr[49469]= 834157373;
assign addr[49470]= 763158411;
assign addr[49471]= 691191324;
assign addr[49472]= 618347408;
assign addr[49473]= 544719071;
assign addr[49474]= 470399716;
assign addr[49475]= 395483624;
assign addr[49476]= 320065829;
assign addr[49477]= 244242007;
assign addr[49478]= 168108346;
assign addr[49479]= 91761426;
assign addr[49480]= 15298099;
assign addr[49481]= -61184634;
assign addr[49482]= -137589750;
assign addr[49483]= -213820322;
assign addr[49484]= -289779648;
assign addr[49485]= -365371365;
assign addr[49486]= -440499581;
assign addr[49487]= -515068990;
assign addr[49488]= -588984994;
assign addr[49489]= -662153826;
assign addr[49490]= -734482665;
assign addr[49491]= -805879757;
assign addr[49492]= -876254528;
assign addr[49493]= -945517704;
assign addr[49494]= -1013581418;
assign addr[49495]= -1080359326;
assign addr[49496]= -1145766716;
assign addr[49497]= -1209720613;
assign addr[49498]= -1272139887;
assign addr[49499]= -1332945355;
assign addr[49500]= -1392059879;
assign addr[49501]= -1449408469;
assign addr[49502]= -1504918373;
assign addr[49503]= -1558519173;
assign addr[49504]= -1610142873;
assign addr[49505]= -1659723983;
assign addr[49506]= -1707199606;
assign addr[49507]= -1752509516;
assign addr[49508]= -1795596234;
assign addr[49509]= -1836405100;
assign addr[49510]= -1874884346;
assign addr[49511]= -1910985158;
assign addr[49512]= -1944661739;
assign addr[49513]= -1975871368;
assign addr[49514]= -2004574453;
assign addr[49515]= -2030734582;
assign addr[49516]= -2054318569;
assign addr[49517]= -2075296495;
assign addr[49518]= -2093641749;
assign addr[49519]= -2109331059;
assign addr[49520]= -2122344521;
assign addr[49521]= -2132665626;
assign addr[49522]= -2140281282;
assign addr[49523]= -2145181827;
assign addr[49524]= -2147361045;
assign addr[49525]= -2146816171;
assign addr[49526]= -2143547897;
assign addr[49527]= -2137560369;
assign addr[49528]= -2128861181;
assign addr[49529]= -2117461370;
assign addr[49530]= -2103375398;
assign addr[49531]= -2086621133;
assign addr[49532]= -2067219829;
assign addr[49533]= -2045196100;
assign addr[49534]= -2020577882;
assign addr[49535]= -1993396407;
assign addr[49536]= -1963686155;
assign addr[49537]= -1931484818;
assign addr[49538]= -1896833245;
assign addr[49539]= -1859775393;
assign addr[49540]= -1820358275;
assign addr[49541]= -1778631892;
assign addr[49542]= -1734649179;
assign addr[49543]= -1688465931;
assign addr[49544]= -1640140734;
assign addr[49545]= -1589734894;
assign addr[49546]= -1537312353;
assign addr[49547]= -1482939614;
assign addr[49548]= -1426685652;
assign addr[49549]= -1368621831;
assign addr[49550]= -1308821808;
assign addr[49551]= -1247361445;
assign addr[49552]= -1184318708;
assign addr[49553]= -1119773573;
assign addr[49554]= -1053807919;
assign addr[49555]= -986505429;
assign addr[49556]= -917951481;
assign addr[49557]= -848233042;
assign addr[49558]= -777438554;
assign addr[49559]= -705657826;
assign addr[49560]= -632981917;
assign addr[49561]= -559503022;
assign addr[49562]= -485314355;
assign addr[49563]= -410510029;
assign addr[49564]= -335184940;
assign addr[49565]= -259434643;
assign addr[49566]= -183355234;
assign addr[49567]= -107043224;
assign addr[49568]= -30595422;
assign addr[49569]= 45891193;
assign addr[49570]= 122319591;
assign addr[49571]= 198592817;
assign addr[49572]= 274614114;
assign addr[49573]= 350287041;
assign addr[49574]= 425515602;
assign addr[49575]= 500204365;
assign addr[49576]= 574258580;
assign addr[49577]= 647584304;
assign addr[49578]= 720088517;
assign addr[49579]= 791679244;
assign addr[49580]= 862265664;
assign addr[49581]= 931758235;
assign addr[49582]= 1000068799;
assign addr[49583]= 1067110699;
assign addr[49584]= 1132798888;
assign addr[49585]= 1197050035;
assign addr[49586]= 1259782632;
assign addr[49587]= 1320917099;
assign addr[49588]= 1380375881;
assign addr[49589]= 1438083551;
assign addr[49590]= 1493966902;
assign addr[49591]= 1547955041;
assign addr[49592]= 1599979481;
assign addr[49593]= 1649974225;
assign addr[49594]= 1697875851;
assign addr[49595]= 1743623590;
assign addr[49596]= 1787159411;
assign addr[49597]= 1828428082;
assign addr[49598]= 1867377253;
assign addr[49599]= 1903957513;
assign addr[49600]= 1938122457;
assign addr[49601]= 1969828744;
assign addr[49602]= 1999036154;
assign addr[49603]= 2025707632;
assign addr[49604]= 2049809346;
assign addr[49605]= 2071310720;
assign addr[49606]= 2090184478;
assign addr[49607]= 2106406677;
assign addr[49608]= 2119956737;
assign addr[49609]= 2130817471;
assign addr[49610]= 2138975100;
assign addr[49611]= 2144419275;
assign addr[49612]= 2147143090;
assign addr[49613]= 2147143090;
assign addr[49614]= 2144419275;
assign addr[49615]= 2138975100;
assign addr[49616]= 2130817471;
assign addr[49617]= 2119956737;
assign addr[49618]= 2106406677;
assign addr[49619]= 2090184478;
assign addr[49620]= 2071310720;
assign addr[49621]= 2049809346;
assign addr[49622]= 2025707632;
assign addr[49623]= 1999036154;
assign addr[49624]= 1969828744;
assign addr[49625]= 1938122457;
assign addr[49626]= 1903957513;
assign addr[49627]= 1867377253;
assign addr[49628]= 1828428082;
assign addr[49629]= 1787159411;
assign addr[49630]= 1743623590;
assign addr[49631]= 1697875851;
assign addr[49632]= 1649974225;
assign addr[49633]= 1599979481;
assign addr[49634]= 1547955041;
assign addr[49635]= 1493966902;
assign addr[49636]= 1438083551;
assign addr[49637]= 1380375881;
assign addr[49638]= 1320917099;
assign addr[49639]= 1259782632;
assign addr[49640]= 1197050035;
assign addr[49641]= 1132798888;
assign addr[49642]= 1067110699;
assign addr[49643]= 1000068799;
assign addr[49644]= 931758235;
assign addr[49645]= 862265664;
assign addr[49646]= 791679244;
assign addr[49647]= 720088517;
assign addr[49648]= 647584304;
assign addr[49649]= 574258580;
assign addr[49650]= 500204365;
assign addr[49651]= 425515602;
assign addr[49652]= 350287041;
assign addr[49653]= 274614114;
assign addr[49654]= 198592817;
assign addr[49655]= 122319591;
assign addr[49656]= 45891193;
assign addr[49657]= -30595422;
assign addr[49658]= -107043224;
assign addr[49659]= -183355234;
assign addr[49660]= -259434643;
assign addr[49661]= -335184940;
assign addr[49662]= -410510029;
assign addr[49663]= -485314355;
assign addr[49664]= -559503022;
assign addr[49665]= -632981917;
assign addr[49666]= -705657826;
assign addr[49667]= -777438554;
assign addr[49668]= -848233042;
assign addr[49669]= -917951481;
assign addr[49670]= -986505429;
assign addr[49671]= -1053807919;
assign addr[49672]= -1119773573;
assign addr[49673]= -1184318708;
assign addr[49674]= -1247361445;
assign addr[49675]= -1308821808;
assign addr[49676]= -1368621831;
assign addr[49677]= -1426685652;
assign addr[49678]= -1482939614;
assign addr[49679]= -1537312353;
assign addr[49680]= -1589734894;
assign addr[49681]= -1640140734;
assign addr[49682]= -1688465931;
assign addr[49683]= -1734649179;
assign addr[49684]= -1778631892;
assign addr[49685]= -1820358275;
assign addr[49686]= -1859775393;
assign addr[49687]= -1896833245;
assign addr[49688]= -1931484818;
assign addr[49689]= -1963686155;
assign addr[49690]= -1993396407;
assign addr[49691]= -2020577882;
assign addr[49692]= -2045196100;
assign addr[49693]= -2067219829;
assign addr[49694]= -2086621133;
assign addr[49695]= -2103375398;
assign addr[49696]= -2117461370;
assign addr[49697]= -2128861181;
assign addr[49698]= -2137560369;
assign addr[49699]= -2143547897;
assign addr[49700]= -2146816171;
assign addr[49701]= -2147361045;
assign addr[49702]= -2145181827;
assign addr[49703]= -2140281282;
assign addr[49704]= -2132665626;
assign addr[49705]= -2122344521;
assign addr[49706]= -2109331059;
assign addr[49707]= -2093641749;
assign addr[49708]= -2075296495;
assign addr[49709]= -2054318569;
assign addr[49710]= -2030734582;
assign addr[49711]= -2004574453;
assign addr[49712]= -1975871368;
assign addr[49713]= -1944661739;
assign addr[49714]= -1910985158;
assign addr[49715]= -1874884346;
assign addr[49716]= -1836405100;
assign addr[49717]= -1795596234;
assign addr[49718]= -1752509516;
assign addr[49719]= -1707199606;
assign addr[49720]= -1659723983;
assign addr[49721]= -1610142873;
assign addr[49722]= -1558519173;
assign addr[49723]= -1504918373;
assign addr[49724]= -1449408469;
assign addr[49725]= -1392059879;
assign addr[49726]= -1332945355;
assign addr[49727]= -1272139887;
assign addr[49728]= -1209720613;
assign addr[49729]= -1145766716;
assign addr[49730]= -1080359326;
assign addr[49731]= -1013581418;
assign addr[49732]= -945517704;
assign addr[49733]= -876254528;
assign addr[49734]= -805879757;
assign addr[49735]= -734482665;
assign addr[49736]= -662153826;
assign addr[49737]= -588984994;
assign addr[49738]= -515068990;
assign addr[49739]= -440499581;
assign addr[49740]= -365371365;
assign addr[49741]= -289779648;
assign addr[49742]= -213820322;
assign addr[49743]= -137589750;
assign addr[49744]= -61184634;
assign addr[49745]= 15298099;
assign addr[49746]= 91761426;
assign addr[49747]= 168108346;
assign addr[49748]= 244242007;
assign addr[49749]= 320065829;
assign addr[49750]= 395483624;
assign addr[49751]= 470399716;
assign addr[49752]= 544719071;
assign addr[49753]= 618347408;
assign addr[49754]= 691191324;
assign addr[49755]= 763158411;
assign addr[49756]= 834157373;
assign addr[49757]= 904098143;
assign addr[49758]= 972891995;
assign addr[49759]= 1040451659;
assign addr[49760]= 1106691431;
assign addr[49761]= 1171527280;
assign addr[49762]= 1234876957;
assign addr[49763]= 1296660098;
assign addr[49764]= 1356798326;
assign addr[49765]= 1415215352;
assign addr[49766]= 1471837070;
assign addr[49767]= 1526591649;
assign addr[49768]= 1579409630;
assign addr[49769]= 1630224009;
assign addr[49770]= 1678970324;
assign addr[49771]= 1725586737;
assign addr[49772]= 1770014111;
assign addr[49773]= 1812196087;
assign addr[49774]= 1852079154;
assign addr[49775]= 1889612716;
assign addr[49776]= 1924749160;
assign addr[49777]= 1957443913;
assign addr[49778]= 1987655498;
assign addr[49779]= 2015345591;
assign addr[49780]= 2040479063;
assign addr[49781]= 2063024031;
assign addr[49782]= 2082951896;
assign addr[49783]= 2100237377;
assign addr[49784]= 2114858546;
assign addr[49785]= 2126796855;
assign addr[49786]= 2136037160;
assign addr[49787]= 2142567738;
assign addr[49788]= 2146380306;
assign addr[49789]= 2147470025;
assign addr[49790]= 2145835515;
assign addr[49791]= 2141478848;
assign addr[49792]= 2134405552;
assign addr[49793]= 2124624598;
assign addr[49794]= 2112148396;
assign addr[49795]= 2096992772;
assign addr[49796]= 2079176953;
assign addr[49797]= 2058723538;
assign addr[49798]= 2035658475;
assign addr[49799]= 2010011024;
assign addr[49800]= 1981813720;
assign addr[49801]= 1951102334;
assign addr[49802]= 1917915825;
assign addr[49803]= 1882296293;
assign addr[49804]= 1844288924;
assign addr[49805]= 1803941934;
assign addr[49806]= 1761306505;
assign addr[49807]= 1716436725;
assign addr[49808]= 1669389513;
assign addr[49809]= 1620224553;
assign addr[49810]= 1569004214;
assign addr[49811]= 1515793473;
assign addr[49812]= 1460659832;
assign addr[49813]= 1403673233;
assign addr[49814]= 1344905966;
assign addr[49815]= 1284432584;
assign addr[49816]= 1222329801;
assign addr[49817]= 1158676398;
assign addr[49818]= 1093553126;
assign addr[49819]= 1027042599;
assign addr[49820]= 959229189;
assign addr[49821]= 890198924;
assign addr[49822]= 820039373;
assign addr[49823]= 748839539;
assign addr[49824]= 676689746;
assign addr[49825]= 603681519;
assign addr[49826]= 529907477;
assign addr[49827]= 455461206;
assign addr[49828]= 380437148;
assign addr[49829]= 304930476;
assign addr[49830]= 229036977;
assign addr[49831]= 152852926;
assign addr[49832]= 76474970;
assign addr[49833]= 0;
assign addr[49834]= -76474970;
assign addr[49835]= -152852926;
assign addr[49836]= -229036977;
assign addr[49837]= -304930476;
assign addr[49838]= -380437148;
assign addr[49839]= -455461206;
assign addr[49840]= -529907477;
assign addr[49841]= -603681519;
assign addr[49842]= -676689746;
assign addr[49843]= -748839539;
assign addr[49844]= -820039373;
assign addr[49845]= -890198924;
assign addr[49846]= -959229189;
assign addr[49847]= -1027042599;
assign addr[49848]= -1093553126;
assign addr[49849]= -1158676398;
assign addr[49850]= -1222329801;
assign addr[49851]= -1284432584;
assign addr[49852]= -1344905966;
assign addr[49853]= -1403673233;
assign addr[49854]= -1460659832;
assign addr[49855]= -1515793473;
assign addr[49856]= -1569004214;
assign addr[49857]= -1620224553;
assign addr[49858]= -1669389513;
assign addr[49859]= -1716436725;
assign addr[49860]= -1761306505;
assign addr[49861]= -1803941934;
assign addr[49862]= -1844288924;
assign addr[49863]= -1882296293;
assign addr[49864]= -1917915825;
assign addr[49865]= -1951102334;
assign addr[49866]= -1981813720;
assign addr[49867]= -2010011024;
assign addr[49868]= -2035658475;
assign addr[49869]= -2058723538;
assign addr[49870]= -2079176953;
assign addr[49871]= -2096992772;
assign addr[49872]= -2112148396;
assign addr[49873]= -2124624598;
assign addr[49874]= -2134405552;
assign addr[49875]= -2141478848;
assign addr[49876]= -2145835515;
assign addr[49877]= -2147470025;
assign addr[49878]= -2146380306;
assign addr[49879]= -2142567738;
assign addr[49880]= -2136037160;
assign addr[49881]= -2126796855;
assign addr[49882]= -2114858546;
assign addr[49883]= -2100237377;
assign addr[49884]= -2082951896;
assign addr[49885]= -2063024031;
assign addr[49886]= -2040479063;
assign addr[49887]= -2015345591;
assign addr[49888]= -1987655498;
assign addr[49889]= -1957443913;
assign addr[49890]= -1924749160;
assign addr[49891]= -1889612716;
assign addr[49892]= -1852079154;
assign addr[49893]= -1812196087;
assign addr[49894]= -1770014111;
assign addr[49895]= -1725586737;
assign addr[49896]= -1678970324;
assign addr[49897]= -1630224009;
assign addr[49898]= -1579409630;
assign addr[49899]= -1526591649;
assign addr[49900]= -1471837070;
assign addr[49901]= -1415215352;
assign addr[49902]= -1356798326;
assign addr[49903]= -1296660098;
assign addr[49904]= -1234876957;
assign addr[49905]= -1171527280;
assign addr[49906]= -1106691431;
assign addr[49907]= -1040451659;
assign addr[49908]= -972891995;
assign addr[49909]= -904098143;
assign addr[49910]= -834157373;
assign addr[49911]= -763158411;
assign addr[49912]= -691191324;
assign addr[49913]= -618347408;
assign addr[49914]= -544719071;
assign addr[49915]= -470399716;
assign addr[49916]= -395483624;
assign addr[49917]= -320065829;
assign addr[49918]= -244242007;
assign addr[49919]= -168108346;
assign addr[49920]= -91761426;
assign addr[49921]= -15298099;
assign addr[49922]= 61184634;
assign addr[49923]= 137589750;
assign addr[49924]= 213820322;
assign addr[49925]= 289779648;
assign addr[49926]= 365371365;
assign addr[49927]= 440499581;
assign addr[49928]= 515068990;
assign addr[49929]= 588984994;
assign addr[49930]= 662153826;
assign addr[49931]= 734482665;
assign addr[49932]= 805879757;
assign addr[49933]= 876254528;
assign addr[49934]= 945517704;
assign addr[49935]= 1013581418;
assign addr[49936]= 1080359326;
assign addr[49937]= 1145766716;
assign addr[49938]= 1209720613;
assign addr[49939]= 1272139887;
assign addr[49940]= 1332945355;
assign addr[49941]= 1392059879;
assign addr[49942]= 1449408469;
assign addr[49943]= 1504918373;
assign addr[49944]= 1558519173;
assign addr[49945]= 1610142873;
assign addr[49946]= 1659723983;
assign addr[49947]= 1707199606;
assign addr[49948]= 1752509516;
assign addr[49949]= 1795596234;
assign addr[49950]= 1836405100;
assign addr[49951]= 1874884346;
assign addr[49952]= 1910985158;
assign addr[49953]= 1944661739;
assign addr[49954]= 1975871368;
assign addr[49955]= 2004574453;
assign addr[49956]= 2030734582;
assign addr[49957]= 2054318569;
assign addr[49958]= 2075296495;
assign addr[49959]= 2093641749;
assign addr[49960]= 2109331059;
assign addr[49961]= 2122344521;
assign addr[49962]= 2132665626;
assign addr[49963]= 2140281282;
assign addr[49964]= 2145181827;
assign addr[49965]= 2147361045;
assign addr[49966]= 2146816171;
assign addr[49967]= 2143547897;
assign addr[49968]= 2137560369;
assign addr[49969]= 2128861181;
assign addr[49970]= 2117461370;
assign addr[49971]= 2103375398;
assign addr[49972]= 2086621133;
assign addr[49973]= 2067219829;
assign addr[49974]= 2045196100;
assign addr[49975]= 2020577882;
assign addr[49976]= 1993396407;
assign addr[49977]= 1963686155;
assign addr[49978]= 1931484818;
assign addr[49979]= 1896833245;
assign addr[49980]= 1859775393;
assign addr[49981]= 1820358275;
assign addr[49982]= 1778631892;
assign addr[49983]= 1734649179;
assign addr[49984]= 1688465931;
assign addr[49985]= 1640140734;
assign addr[49986]= 1589734894;
assign addr[49987]= 1537312353;
assign addr[49988]= 1482939614;
assign addr[49989]= 1426685652;
assign addr[49990]= 1368621831;
assign addr[49991]= 1308821808;
assign addr[49992]= 1247361445;
assign addr[49993]= 1184318708;
assign addr[49994]= 1119773573;
assign addr[49995]= 1053807919;
assign addr[49996]= 986505429;
assign addr[49997]= 917951481;
assign addr[49998]= 848233042;
assign addr[49999]= 777438554;
assign addr[50000]= 705657826;
assign addr[50001]= 632981917;
assign addr[50002]= 559503022;
assign addr[50003]= 485314355;
assign addr[50004]= 410510029;
assign addr[50005]= 335184940;
assign addr[50006]= 259434643;
assign addr[50007]= 183355234;
assign addr[50008]= 107043224;
assign addr[50009]= 30595422;
assign addr[50010]= -45891193;
assign addr[50011]= -122319591;
assign addr[50012]= -198592817;
assign addr[50013]= -274614114;
assign addr[50014]= -350287041;
assign addr[50015]= -425515602;
assign addr[50016]= -500204365;
assign addr[50017]= -574258580;
assign addr[50018]= -647584304;
assign addr[50019]= -720088517;
assign addr[50020]= -791679244;
assign addr[50021]= -862265664;
assign addr[50022]= -931758235;
assign addr[50023]= -1000068799;
assign addr[50024]= -1067110699;
assign addr[50025]= -1132798888;
assign addr[50026]= -1197050035;
assign addr[50027]= -1259782632;
assign addr[50028]= -1320917099;
assign addr[50029]= -1380375881;
assign addr[50030]= -1438083551;
assign addr[50031]= -1493966902;
assign addr[50032]= -1547955041;
assign addr[50033]= -1599979481;
assign addr[50034]= -1649974225;
assign addr[50035]= -1697875851;
assign addr[50036]= -1743623590;
assign addr[50037]= -1787159411;
assign addr[50038]= -1828428082;
assign addr[50039]= -1867377253;
assign addr[50040]= -1903957513;
assign addr[50041]= -1938122457;
assign addr[50042]= -1969828744;
assign addr[50043]= -1999036154;
assign addr[50044]= -2025707632;
assign addr[50045]= -2049809346;
assign addr[50046]= -2071310720;
assign addr[50047]= -2090184478;
assign addr[50048]= -2106406677;
assign addr[50049]= -2119956737;
assign addr[50050]= -2130817471;
assign addr[50051]= -2138975100;
assign addr[50052]= -2144419275;
assign addr[50053]= -2147143090;
assign addr[50054]= -2147143090;
assign addr[50055]= -2144419275;
assign addr[50056]= -2138975100;
assign addr[50057]= -2130817471;
assign addr[50058]= -2119956737;
assign addr[50059]= -2106406677;
assign addr[50060]= -2090184478;
assign addr[50061]= -2071310720;
assign addr[50062]= -2049809346;
assign addr[50063]= -2025707632;
assign addr[50064]= -1999036154;
assign addr[50065]= -1969828744;
assign addr[50066]= -1938122457;
assign addr[50067]= -1903957513;
assign addr[50068]= -1867377253;
assign addr[50069]= -1828428082;
assign addr[50070]= -1787159411;
assign addr[50071]= -1743623590;
assign addr[50072]= -1697875851;
assign addr[50073]= -1649974225;
assign addr[50074]= -1599979481;
assign addr[50075]= -1547955041;
assign addr[50076]= -1493966902;
assign addr[50077]= -1438083551;
assign addr[50078]= -1380375881;
assign addr[50079]= -1320917099;
assign addr[50080]= -1259782632;
assign addr[50081]= -1197050035;
assign addr[50082]= -1132798888;
assign addr[50083]= -1067110699;
assign addr[50084]= -1000068799;
assign addr[50085]= -931758235;
assign addr[50086]= -862265664;
assign addr[50087]= -791679244;
assign addr[50088]= -720088517;
assign addr[50089]= -647584304;
assign addr[50090]= -574258580;
assign addr[50091]= -500204365;
assign addr[50092]= -425515602;
assign addr[50093]= -350287041;
assign addr[50094]= -274614114;
assign addr[50095]= -198592817;
assign addr[50096]= -122319591;
assign addr[50097]= -45891193;
assign addr[50098]= 30595422;
assign addr[50099]= 107043224;
assign addr[50100]= 183355234;
assign addr[50101]= 259434643;
assign addr[50102]= 335184940;
assign addr[50103]= 410510029;
assign addr[50104]= 485314355;
assign addr[50105]= 559503022;
assign addr[50106]= 632981917;
assign addr[50107]= 705657826;
assign addr[50108]= 777438554;
assign addr[50109]= 848233042;
assign addr[50110]= 917951481;
assign addr[50111]= 986505429;
assign addr[50112]= 1053807919;
assign addr[50113]= 1119773573;
assign addr[50114]= 1184318708;
assign addr[50115]= 1247361445;
assign addr[50116]= 1308821808;
assign addr[50117]= 1368621831;
assign addr[50118]= 1426685652;
assign addr[50119]= 1482939614;
assign addr[50120]= 1537312353;
assign addr[50121]= 1589734894;
assign addr[50122]= 1640140734;
assign addr[50123]= 1688465931;
assign addr[50124]= 1734649179;
assign addr[50125]= 1778631892;
assign addr[50126]= 1820358275;
assign addr[50127]= 1859775393;
assign addr[50128]= 1896833245;
assign addr[50129]= 1931484818;
assign addr[50130]= 1963686155;
assign addr[50131]= 1993396407;
assign addr[50132]= 2020577882;
assign addr[50133]= 2045196100;
assign addr[50134]= 2067219829;
assign addr[50135]= 2086621133;
assign addr[50136]= 2103375398;
assign addr[50137]= 2117461370;
assign addr[50138]= 2128861181;
assign addr[50139]= 2137560369;
assign addr[50140]= 2143547897;
assign addr[50141]= 2146816171;
assign addr[50142]= 2147361045;
assign addr[50143]= 2145181827;
assign addr[50144]= 2140281282;
assign addr[50145]= 2132665626;
assign addr[50146]= 2122344521;
assign addr[50147]= 2109331059;
assign addr[50148]= 2093641749;
assign addr[50149]= 2075296495;
assign addr[50150]= 2054318569;
assign addr[50151]= 2030734582;
assign addr[50152]= 2004574453;
assign addr[50153]= 1975871368;
assign addr[50154]= 1944661739;
assign addr[50155]= 1910985158;
assign addr[50156]= 1874884346;
assign addr[50157]= 1836405100;
assign addr[50158]= 1795596234;
assign addr[50159]= 1752509516;
assign addr[50160]= 1707199606;
assign addr[50161]= 1659723983;
assign addr[50162]= 1610142873;
assign addr[50163]= 1558519173;
assign addr[50164]= 1504918373;
assign addr[50165]= 1449408469;
assign addr[50166]= 1392059879;
assign addr[50167]= 1332945355;
assign addr[50168]= 1272139887;
assign addr[50169]= 1209720613;
assign addr[50170]= 1145766716;
assign addr[50171]= 1080359326;
assign addr[50172]= 1013581418;
assign addr[50173]= 945517704;
assign addr[50174]= 876254528;
assign addr[50175]= 805879757;
assign addr[50176]= 734482665;
assign addr[50177]= 662153826;
assign addr[50178]= 588984994;
assign addr[50179]= 515068990;
assign addr[50180]= 440499581;
assign addr[50181]= 365371365;
assign addr[50182]= 289779648;
assign addr[50183]= 213820322;
assign addr[50184]= 137589750;
assign addr[50185]= 61184634;
assign addr[50186]= -15298099;
assign addr[50187]= -91761426;
assign addr[50188]= -168108346;
assign addr[50189]= -244242007;
assign addr[50190]= -320065829;
assign addr[50191]= -395483624;
assign addr[50192]= -470399716;
assign addr[50193]= -544719071;
assign addr[50194]= -618347408;
assign addr[50195]= -691191324;
assign addr[50196]= -763158411;
assign addr[50197]= -834157373;
assign addr[50198]= -904098143;
assign addr[50199]= -972891995;
assign addr[50200]= -1040451659;
assign addr[50201]= -1106691431;
assign addr[50202]= -1171527280;
assign addr[50203]= -1234876957;
assign addr[50204]= -1296660098;
assign addr[50205]= -1356798326;
assign addr[50206]= -1415215352;
assign addr[50207]= -1471837070;
assign addr[50208]= -1526591649;
assign addr[50209]= -1579409630;
assign addr[50210]= -1630224009;
assign addr[50211]= -1678970324;
assign addr[50212]= -1725586737;
assign addr[50213]= -1770014111;
assign addr[50214]= -1812196087;
assign addr[50215]= -1852079154;
assign addr[50216]= -1889612716;
assign addr[50217]= -1924749160;
assign addr[50218]= -1957443913;
assign addr[50219]= -1987655498;
assign addr[50220]= -2015345591;
assign addr[50221]= -2040479063;
assign addr[50222]= -2063024031;
assign addr[50223]= -2082951896;
assign addr[50224]= -2100237377;
assign addr[50225]= -2114858546;
assign addr[50226]= -2126796855;
assign addr[50227]= -2136037160;
assign addr[50228]= -2142567738;
assign addr[50229]= -2146380306;
assign addr[50230]= -2147470025;
assign addr[50231]= -2145835515;
assign addr[50232]= -2141478848;
assign addr[50233]= -2134405552;
assign addr[50234]= -2124624598;
assign addr[50235]= -2112148396;
assign addr[50236]= -2096992772;
assign addr[50237]= -2079176953;
assign addr[50238]= -2058723538;
assign addr[50239]= -2035658475;
assign addr[50240]= -2010011024;
assign addr[50241]= -1981813720;
assign addr[50242]= -1951102334;
assign addr[50243]= -1917915825;
assign addr[50244]= -1882296293;
assign addr[50245]= -1844288924;
assign addr[50246]= -1803941934;
assign addr[50247]= -1761306505;
assign addr[50248]= -1716436725;
assign addr[50249]= -1669389513;
assign addr[50250]= -1620224553;
assign addr[50251]= -1569004214;
assign addr[50252]= -1515793473;
assign addr[50253]= -1460659832;
assign addr[50254]= -1403673233;
assign addr[50255]= -1344905966;
assign addr[50256]= -1284432584;
assign addr[50257]= -1222329801;
assign addr[50258]= -1158676398;
assign addr[50259]= -1093553126;
assign addr[50260]= -1027042599;
assign addr[50261]= -959229189;
assign addr[50262]= -890198924;
assign addr[50263]= -820039373;
assign addr[50264]= -748839539;
assign addr[50265]= -676689746;
assign addr[50266]= -603681519;
assign addr[50267]= -529907477;
assign addr[50268]= -455461206;
assign addr[50269]= -380437148;
assign addr[50270]= -304930476;
assign addr[50271]= -229036977;
assign addr[50272]= -152852926;
assign addr[50273]= -76474970;
assign addr[50274]= 0;
assign addr[50275]= 76474970;
assign addr[50276]= 152852926;
assign addr[50277]= 229036977;
assign addr[50278]= 304930476;
assign addr[50279]= 380437148;
assign addr[50280]= 455461206;
assign addr[50281]= 529907477;
assign addr[50282]= 603681519;
assign addr[50283]= 676689746;
assign addr[50284]= 748839539;
assign addr[50285]= 820039373;
assign addr[50286]= 890198924;
assign addr[50287]= 959229189;
assign addr[50288]= 1027042599;
assign addr[50289]= 1093553126;
assign addr[50290]= 1158676398;
assign addr[50291]= 1222329801;
assign addr[50292]= 1284432584;
assign addr[50293]= 1344905966;
assign addr[50294]= 1403673233;
assign addr[50295]= 1460659832;
assign addr[50296]= 1515793473;
assign addr[50297]= 1569004214;
assign addr[50298]= 1620224553;
assign addr[50299]= 1669389513;
assign addr[50300]= 1716436725;
assign addr[50301]= 1761306505;
assign addr[50302]= 1803941934;
assign addr[50303]= 1844288924;
assign addr[50304]= 1882296293;
assign addr[50305]= 1917915825;
assign addr[50306]= 1951102334;
assign addr[50307]= 1981813720;
assign addr[50308]= 2010011024;
assign addr[50309]= 2035658475;
assign addr[50310]= 2058723538;
assign addr[50311]= 2079176953;
assign addr[50312]= 2096992772;
assign addr[50313]= 2112148396;
assign addr[50314]= 2124624598;
assign addr[50315]= 2134405552;
assign addr[50316]= 2141478848;
assign addr[50317]= 2145835515;
assign addr[50318]= 2147470025;
assign addr[50319]= 2146380306;
assign addr[50320]= 2142567738;
assign addr[50321]= 2136037160;
assign addr[50322]= 2126796855;
assign addr[50323]= 2114858546;
assign addr[50324]= 2100237377;
assign addr[50325]= 2082951896;
assign addr[50326]= 2063024031;
assign addr[50327]= 2040479063;
assign addr[50328]= 2015345591;
assign addr[50329]= 1987655498;
assign addr[50330]= 1957443913;
assign addr[50331]= 1924749160;
assign addr[50332]= 1889612716;
assign addr[50333]= 1852079154;
assign addr[50334]= 1812196087;
assign addr[50335]= 1770014111;
assign addr[50336]= 1725586737;
assign addr[50337]= 1678970324;
assign addr[50338]= 1630224009;
assign addr[50339]= 1579409630;
assign addr[50340]= 1526591649;
assign addr[50341]= 1471837070;
assign addr[50342]= 1415215352;
assign addr[50343]= 1356798326;
assign addr[50344]= 1296660098;
assign addr[50345]= 1234876957;
assign addr[50346]= 1171527280;
assign addr[50347]= 1106691431;
assign addr[50348]= 1040451659;
assign addr[50349]= 972891995;
assign addr[50350]= 904098143;
assign addr[50351]= 834157373;
assign addr[50352]= 763158411;
assign addr[50353]= 691191324;
assign addr[50354]= 618347408;
assign addr[50355]= 544719071;
assign addr[50356]= 470399716;
assign addr[50357]= 395483624;
assign addr[50358]= 320065829;
assign addr[50359]= 244242007;
assign addr[50360]= 168108346;
assign addr[50361]= 91761426;
assign addr[50362]= 15298099;
assign addr[50363]= -61184634;
assign addr[50364]= -137589750;
assign addr[50365]= -213820322;
assign addr[50366]= -289779648;
assign addr[50367]= -365371365;
assign addr[50368]= -440499581;
assign addr[50369]= -515068990;
assign addr[50370]= -588984994;
assign addr[50371]= -662153826;
assign addr[50372]= -734482665;
assign addr[50373]= -805879757;
assign addr[50374]= -876254528;
assign addr[50375]= -945517704;
assign addr[50376]= -1013581418;
assign addr[50377]= -1080359326;
assign addr[50378]= -1145766716;
assign addr[50379]= -1209720613;
assign addr[50380]= -1272139887;
assign addr[50381]= -1332945355;
assign addr[50382]= -1392059879;
assign addr[50383]= -1449408469;
assign addr[50384]= -1504918373;
assign addr[50385]= -1558519173;
assign addr[50386]= -1610142873;
assign addr[50387]= -1659723983;
assign addr[50388]= -1707199606;
assign addr[50389]= -1752509516;
assign addr[50390]= -1795596234;
assign addr[50391]= -1836405100;
assign addr[50392]= -1874884346;
assign addr[50393]= -1910985158;
assign addr[50394]= -1944661739;
assign addr[50395]= -1975871368;
assign addr[50396]= -2004574453;
assign addr[50397]= -2030734582;
assign addr[50398]= -2054318569;
assign addr[50399]= -2075296495;
assign addr[50400]= -2093641749;
assign addr[50401]= -2109331059;
assign addr[50402]= -2122344521;
assign addr[50403]= -2132665626;
assign addr[50404]= -2140281282;
assign addr[50405]= -2145181827;
assign addr[50406]= -2147361045;
assign addr[50407]= -2146816171;
assign addr[50408]= -2143547897;
assign addr[50409]= -2137560369;
assign addr[50410]= -2128861181;
assign addr[50411]= -2117461370;
assign addr[50412]= -2103375398;
assign addr[50413]= -2086621133;
assign addr[50414]= -2067219829;
assign addr[50415]= -2045196100;
assign addr[50416]= -2020577882;
assign addr[50417]= -1993396407;
assign addr[50418]= -1963686155;
assign addr[50419]= -1931484818;
assign addr[50420]= -1896833245;
assign addr[50421]= -1859775393;
assign addr[50422]= -1820358275;
assign addr[50423]= -1778631892;
assign addr[50424]= -1734649179;
assign addr[50425]= -1688465931;
assign addr[50426]= -1640140734;
assign addr[50427]= -1589734894;
assign addr[50428]= -1537312353;
assign addr[50429]= -1482939614;
assign addr[50430]= -1426685652;
assign addr[50431]= -1368621831;
assign addr[50432]= -1308821808;
assign addr[50433]= -1247361445;
assign addr[50434]= -1184318708;
assign addr[50435]= -1119773573;
assign addr[50436]= -1053807919;
assign addr[50437]= -986505429;
assign addr[50438]= -917951481;
assign addr[50439]= -848233042;
assign addr[50440]= -777438554;
assign addr[50441]= -705657826;
assign addr[50442]= -632981917;
assign addr[50443]= -559503022;
assign addr[50444]= -485314355;
assign addr[50445]= -410510029;
assign addr[50446]= -335184940;
assign addr[50447]= -259434643;
assign addr[50448]= -183355234;
assign addr[50449]= -107043224;
assign addr[50450]= -30595422;
assign addr[50451]= 45891193;
assign addr[50452]= 122319591;
assign addr[50453]= 198592817;
assign addr[50454]= 274614114;
assign addr[50455]= 350287041;
assign addr[50456]= 425515602;
assign addr[50457]= 500204365;
assign addr[50458]= 574258580;
assign addr[50459]= 647584304;
assign addr[50460]= 720088517;
assign addr[50461]= 791679244;
assign addr[50462]= 862265664;
assign addr[50463]= 931758235;
assign addr[50464]= 1000068799;
assign addr[50465]= 1067110699;
assign addr[50466]= 1132798888;
assign addr[50467]= 1197050035;
assign addr[50468]= 1259782632;
assign addr[50469]= 1320917099;
assign addr[50470]= 1380375881;
assign addr[50471]= 1438083551;
assign addr[50472]= 1493966902;
assign addr[50473]= 1547955041;
assign addr[50474]= 1599979481;
assign addr[50475]= 1649974225;
assign addr[50476]= 1697875851;
assign addr[50477]= 1743623590;
assign addr[50478]= 1787159411;
assign addr[50479]= 1828428082;
assign addr[50480]= 1867377253;
assign addr[50481]= 1903957513;
assign addr[50482]= 1938122457;
assign addr[50483]= 1969828744;
assign addr[50484]= 1999036154;
assign addr[50485]= 2025707632;
assign addr[50486]= 2049809346;
assign addr[50487]= 2071310720;
assign addr[50488]= 2090184478;
assign addr[50489]= 2106406677;
assign addr[50490]= 2119956737;
assign addr[50491]= 2130817471;
assign addr[50492]= 2138975100;
assign addr[50493]= 2144419275;
assign addr[50494]= 2147143090;
assign addr[50495]= 2147143090;
assign addr[50496]= 2144419275;
assign addr[50497]= 2138975100;
assign addr[50498]= 2130817471;
assign addr[50499]= 2119956737;
assign addr[50500]= 2106406677;
assign addr[50501]= 2090184478;
assign addr[50502]= 2071310720;
assign addr[50503]= 2049809346;
assign addr[50504]= 2025707632;
assign addr[50505]= 1999036154;
assign addr[50506]= 1969828744;
assign addr[50507]= 1938122457;
assign addr[50508]= 1903957513;
assign addr[50509]= 1867377253;
assign addr[50510]= 1828428082;
assign addr[50511]= 1787159411;
assign addr[50512]= 1743623590;
assign addr[50513]= 1697875851;
assign addr[50514]= 1649974225;
assign addr[50515]= 1599979481;
assign addr[50516]= 1547955041;
assign addr[50517]= 1493966902;
assign addr[50518]= 1438083551;
assign addr[50519]= 1380375881;
assign addr[50520]= 1320917099;
assign addr[50521]= 1259782632;
assign addr[50522]= 1197050035;
assign addr[50523]= 1132798888;
assign addr[50524]= 1067110699;
assign addr[50525]= 1000068799;
assign addr[50526]= 931758235;
assign addr[50527]= 862265664;
assign addr[50528]= 791679244;
assign addr[50529]= 720088517;
assign addr[50530]= 647584304;
assign addr[50531]= 574258580;
assign addr[50532]= 500204365;
assign addr[50533]= 425515602;
assign addr[50534]= 350287041;
assign addr[50535]= 274614114;
assign addr[50536]= 198592817;
assign addr[50537]= 122319591;
assign addr[50538]= 45891193;
assign addr[50539]= -30595422;
assign addr[50540]= -107043224;
assign addr[50541]= -183355234;
assign addr[50542]= -259434643;
assign addr[50543]= -335184940;
assign addr[50544]= -410510029;
assign addr[50545]= -485314355;
assign addr[50546]= -559503022;
assign addr[50547]= -632981917;
assign addr[50548]= -705657826;
assign addr[50549]= -777438554;
assign addr[50550]= -848233042;
assign addr[50551]= -917951481;
assign addr[50552]= -986505429;
assign addr[50553]= -1053807919;
assign addr[50554]= -1119773573;
assign addr[50555]= -1184318708;
assign addr[50556]= -1247361445;
assign addr[50557]= -1308821808;
assign addr[50558]= -1368621831;
assign addr[50559]= -1426685652;
assign addr[50560]= -1482939614;
assign addr[50561]= -1537312353;
assign addr[50562]= -1589734894;
assign addr[50563]= -1640140734;
assign addr[50564]= -1688465931;
assign addr[50565]= -1734649179;
assign addr[50566]= -1778631892;
assign addr[50567]= -1820358275;
assign addr[50568]= -1859775393;
assign addr[50569]= -1896833245;
assign addr[50570]= -1931484818;
assign addr[50571]= -1963686155;
assign addr[50572]= -1993396407;
assign addr[50573]= -2020577882;
assign addr[50574]= -2045196100;
assign addr[50575]= -2067219829;
assign addr[50576]= -2086621133;
assign addr[50577]= -2103375398;
assign addr[50578]= -2117461370;
assign addr[50579]= -2128861181;
assign addr[50580]= -2137560369;
assign addr[50581]= -2143547897;
assign addr[50582]= -2146816171;
assign addr[50583]= -2147361045;
assign addr[50584]= -2145181827;
assign addr[50585]= -2140281282;
assign addr[50586]= -2132665626;
assign addr[50587]= -2122344521;
assign addr[50588]= -2109331059;
assign addr[50589]= -2093641749;
assign addr[50590]= -2075296495;
assign addr[50591]= -2054318569;
assign addr[50592]= -2030734582;
assign addr[50593]= -2004574453;
assign addr[50594]= -1975871368;
assign addr[50595]= -1944661739;
assign addr[50596]= -1910985158;
assign addr[50597]= -1874884346;
assign addr[50598]= -1836405100;
assign addr[50599]= -1795596234;
assign addr[50600]= -1752509516;
assign addr[50601]= -1707199606;
assign addr[50602]= -1659723983;
assign addr[50603]= -1610142873;
assign addr[50604]= -1558519173;
assign addr[50605]= -1504918373;
assign addr[50606]= -1449408469;
assign addr[50607]= -1392059879;
assign addr[50608]= -1332945355;
assign addr[50609]= -1272139887;
assign addr[50610]= -1209720613;
assign addr[50611]= -1145766716;
assign addr[50612]= -1080359326;
assign addr[50613]= -1013581418;
assign addr[50614]= -945517704;
assign addr[50615]= -876254528;
assign addr[50616]= -805879757;
assign addr[50617]= -734482665;
assign addr[50618]= -662153826;
assign addr[50619]= -588984994;
assign addr[50620]= -515068990;
assign addr[50621]= -440499581;
assign addr[50622]= -365371365;
assign addr[50623]= -289779648;
assign addr[50624]= -213820322;
assign addr[50625]= -137589750;
assign addr[50626]= -61184634;
assign addr[50627]= 15298099;
assign addr[50628]= 91761426;
assign addr[50629]= 168108346;
assign addr[50630]= 244242007;
assign addr[50631]= 320065829;
assign addr[50632]= 395483624;
assign addr[50633]= 470399716;
assign addr[50634]= 544719071;
assign addr[50635]= 618347408;
assign addr[50636]= 691191324;
assign addr[50637]= 763158411;
assign addr[50638]= 834157373;
assign addr[50639]= 904098143;
assign addr[50640]= 972891995;
assign addr[50641]= 1040451659;
assign addr[50642]= 1106691431;
assign addr[50643]= 1171527280;
assign addr[50644]= 1234876957;
assign addr[50645]= 1296660098;
assign addr[50646]= 1356798326;
assign addr[50647]= 1415215352;
assign addr[50648]= 1471837070;
assign addr[50649]= 1526591649;
assign addr[50650]= 1579409630;
assign addr[50651]= 1630224009;
assign addr[50652]= 1678970324;
assign addr[50653]= 1725586737;
assign addr[50654]= 1770014111;
assign addr[50655]= 1812196087;
assign addr[50656]= 1852079154;
assign addr[50657]= 1889612716;
assign addr[50658]= 1924749160;
assign addr[50659]= 1957443913;
assign addr[50660]= 1987655498;
assign addr[50661]= 2015345591;
assign addr[50662]= 2040479063;
assign addr[50663]= 2063024031;
assign addr[50664]= 2082951896;
assign addr[50665]= 2100237377;
assign addr[50666]= 2114858546;
assign addr[50667]= 2126796855;
assign addr[50668]= 2136037160;
assign addr[50669]= 2142567738;
assign addr[50670]= 2146380306;
assign addr[50671]= 2147470025;
assign addr[50672]= 2145835515;
assign addr[50673]= 2141478848;
assign addr[50674]= 2134405552;
assign addr[50675]= 2124624598;
assign addr[50676]= 2112148396;
assign addr[50677]= 2096992772;
assign addr[50678]= 2079176953;
assign addr[50679]= 2058723538;
assign addr[50680]= 2035658475;
assign addr[50681]= 2010011024;
assign addr[50682]= 1981813720;
assign addr[50683]= 1951102334;
assign addr[50684]= 1917915825;
assign addr[50685]= 1882296293;
assign addr[50686]= 1844288924;
assign addr[50687]= 1803941934;
assign addr[50688]= 1761306505;
assign addr[50689]= 1716436725;
assign addr[50690]= 1669389513;
assign addr[50691]= 1620224553;
assign addr[50692]= 1569004214;
assign addr[50693]= 1515793473;
assign addr[50694]= 1460659832;
assign addr[50695]= 1403673233;
assign addr[50696]= 1344905966;
assign addr[50697]= 1284432584;
assign addr[50698]= 1222329801;
assign addr[50699]= 1158676398;
assign addr[50700]= 1093553126;
assign addr[50701]= 1027042599;
assign addr[50702]= 959229189;
assign addr[50703]= 890198924;
assign addr[50704]= 820039373;
assign addr[50705]= 748839539;
assign addr[50706]= 676689746;
assign addr[50707]= 603681519;
assign addr[50708]= 529907477;
assign addr[50709]= 455461206;
assign addr[50710]= 380437148;
assign addr[50711]= 304930476;
assign addr[50712]= 229036977;
assign addr[50713]= 152852926;
assign addr[50714]= 76474970;
assign addr[50715]= 0;
assign addr[50716]= -76474970;
assign addr[50717]= -152852926;
assign addr[50718]= -229036977;
assign addr[50719]= -304930476;
assign addr[50720]= -380437148;
assign addr[50721]= -455461206;
assign addr[50722]= -529907477;
assign addr[50723]= -603681519;
assign addr[50724]= -676689746;
assign addr[50725]= -748839539;
assign addr[50726]= -820039373;
assign addr[50727]= -890198924;
assign addr[50728]= -959229189;
assign addr[50729]= -1027042599;
assign addr[50730]= -1093553126;
assign addr[50731]= -1158676398;
assign addr[50732]= -1222329801;
assign addr[50733]= -1284432584;
assign addr[50734]= -1344905966;
assign addr[50735]= -1403673233;
assign addr[50736]= -1460659832;
assign addr[50737]= -1515793473;
assign addr[50738]= -1569004214;
assign addr[50739]= -1620224553;
assign addr[50740]= -1669389513;
assign addr[50741]= -1716436725;
assign addr[50742]= -1761306505;
assign addr[50743]= -1803941934;
assign addr[50744]= -1844288924;
assign addr[50745]= -1882296293;
assign addr[50746]= -1917915825;
assign addr[50747]= -1951102334;
assign addr[50748]= -1981813720;
assign addr[50749]= -2010011024;
assign addr[50750]= -2035658475;
assign addr[50751]= -2058723538;
assign addr[50752]= -2079176953;
assign addr[50753]= -2096992772;
assign addr[50754]= -2112148396;
assign addr[50755]= -2124624598;
assign addr[50756]= -2134405552;
assign addr[50757]= -2141478848;
assign addr[50758]= -2145835515;
assign addr[50759]= -2147470025;
assign addr[50760]= -2146380306;
assign addr[50761]= -2142567738;
assign addr[50762]= -2136037160;
assign addr[50763]= -2126796855;
assign addr[50764]= -2114858546;
assign addr[50765]= -2100237377;
assign addr[50766]= -2082951896;
assign addr[50767]= -2063024031;
assign addr[50768]= -2040479063;
assign addr[50769]= -2015345591;
assign addr[50770]= -1987655498;
assign addr[50771]= -1957443913;
assign addr[50772]= -1924749160;
assign addr[50773]= -1889612716;
assign addr[50774]= -1852079154;
assign addr[50775]= -1812196087;
assign addr[50776]= -1770014111;
assign addr[50777]= -1725586737;
assign addr[50778]= -1678970324;
assign addr[50779]= -1630224009;
assign addr[50780]= -1579409630;
assign addr[50781]= -1526591649;
assign addr[50782]= -1471837070;
assign addr[50783]= -1415215352;
assign addr[50784]= -1356798326;
assign addr[50785]= -1296660098;
assign addr[50786]= -1234876957;
assign addr[50787]= -1171527280;
assign addr[50788]= -1106691431;
assign addr[50789]= -1040451659;
assign addr[50790]= -972891995;
assign addr[50791]= -904098143;
assign addr[50792]= -834157373;
assign addr[50793]= -763158411;
assign addr[50794]= -691191324;
assign addr[50795]= -618347408;
assign addr[50796]= -544719071;
assign addr[50797]= -470399716;
assign addr[50798]= -395483624;
assign addr[50799]= -320065829;
assign addr[50800]= -244242007;
assign addr[50801]= -168108346;
assign addr[50802]= -91761426;
assign addr[50803]= -15298099;
assign addr[50804]= 61184634;
assign addr[50805]= 137589750;
assign addr[50806]= 213820322;
assign addr[50807]= 289779648;
assign addr[50808]= 365371365;
assign addr[50809]= 440499581;
assign addr[50810]= 515068990;
assign addr[50811]= 588984994;
assign addr[50812]= 662153826;
assign addr[50813]= 734482665;
assign addr[50814]= 805879757;
assign addr[50815]= 876254528;
assign addr[50816]= 945517704;
assign addr[50817]= 1013581418;
assign addr[50818]= 1080359326;
assign addr[50819]= 1145766716;
assign addr[50820]= 1209720613;
assign addr[50821]= 1272139887;
assign addr[50822]= 1332945355;
assign addr[50823]= 1392059879;
assign addr[50824]= 1449408469;
assign addr[50825]= 1504918373;
assign addr[50826]= 1558519173;
assign addr[50827]= 1610142873;
assign addr[50828]= 1659723983;
assign addr[50829]= 1707199606;
assign addr[50830]= 1752509516;
assign addr[50831]= 1795596234;
assign addr[50832]= 1836405100;
assign addr[50833]= 1874884346;
assign addr[50834]= 1910985158;
assign addr[50835]= 1944661739;
assign addr[50836]= 1975871368;
assign addr[50837]= 2004574453;
assign addr[50838]= 2030734582;
assign addr[50839]= 2054318569;
assign addr[50840]= 2075296495;
assign addr[50841]= 2093641749;
assign addr[50842]= 2109331059;
assign addr[50843]= 2122344521;
assign addr[50844]= 2132665626;
assign addr[50845]= 2140281282;
assign addr[50846]= 2145181827;
assign addr[50847]= 2147361045;
assign addr[50848]= 2146816171;
assign addr[50849]= 2143547897;
assign addr[50850]= 2137560369;
assign addr[50851]= 2128861181;
assign addr[50852]= 2117461370;
assign addr[50853]= 2103375398;
assign addr[50854]= 2086621133;
assign addr[50855]= 2067219829;
assign addr[50856]= 2045196100;
assign addr[50857]= 2020577882;
assign addr[50858]= 1993396407;
assign addr[50859]= 1963686155;
assign addr[50860]= 1931484818;
assign addr[50861]= 1896833245;
assign addr[50862]= 1859775393;
assign addr[50863]= 1820358275;
assign addr[50864]= 1778631892;
assign addr[50865]= 1734649179;
assign addr[50866]= 1688465931;
assign addr[50867]= 1640140734;
assign addr[50868]= 1589734894;
assign addr[50869]= 1537312353;
assign addr[50870]= 1482939614;
assign addr[50871]= 1426685652;
assign addr[50872]= 1368621831;
assign addr[50873]= 1308821808;
assign addr[50874]= 1247361445;
assign addr[50875]= 1184318708;
assign addr[50876]= 1119773573;
assign addr[50877]= 1053807919;
assign addr[50878]= 986505429;
assign addr[50879]= 917951481;
assign addr[50880]= 848233042;
assign addr[50881]= 777438554;
assign addr[50882]= 705657826;
assign addr[50883]= 632981917;
assign addr[50884]= 559503022;
assign addr[50885]= 485314355;
assign addr[50886]= 410510029;
assign addr[50887]= 335184940;
assign addr[50888]= 259434643;
assign addr[50889]= 183355234;
assign addr[50890]= 107043224;
assign addr[50891]= 30595422;
assign addr[50892]= -45891193;
assign addr[50893]= -122319591;
assign addr[50894]= -198592817;
assign addr[50895]= -274614114;
assign addr[50896]= -350287041;
assign addr[50897]= -425515602;
assign addr[50898]= -500204365;
assign addr[50899]= -574258580;
assign addr[50900]= -647584304;
assign addr[50901]= -720088517;
assign addr[50902]= -791679244;
assign addr[50903]= -862265664;
assign addr[50904]= -931758235;
assign addr[50905]= -1000068799;
assign addr[50906]= -1067110699;
assign addr[50907]= -1132798888;
assign addr[50908]= -1197050035;
assign addr[50909]= -1259782632;
assign addr[50910]= -1320917099;
assign addr[50911]= -1380375881;
assign addr[50912]= -1438083551;
assign addr[50913]= -1493966902;
assign addr[50914]= -1547955041;
assign addr[50915]= -1599979481;
assign addr[50916]= -1649974225;
assign addr[50917]= -1697875851;
assign addr[50918]= -1743623590;
assign addr[50919]= -1787159411;
assign addr[50920]= -1828428082;
assign addr[50921]= -1867377253;
assign addr[50922]= -1903957513;
assign addr[50923]= -1938122457;
assign addr[50924]= -1969828744;
assign addr[50925]= -1999036154;
assign addr[50926]= -2025707632;
assign addr[50927]= -2049809346;
assign addr[50928]= -2071310720;
assign addr[50929]= -2090184478;
assign addr[50930]= -2106406677;
assign addr[50931]= -2119956737;
assign addr[50932]= -2130817471;
assign addr[50933]= -2138975100;
assign addr[50934]= -2144419275;
assign addr[50935]= -2147143090;
assign addr[50936]= -2147143090;
assign addr[50937]= -2144419275;
assign addr[50938]= -2138975100;
assign addr[50939]= -2130817471;
assign addr[50940]= -2119956737;
assign addr[50941]= -2106406677;
assign addr[50942]= -2090184478;
assign addr[50943]= -2071310720;
assign addr[50944]= -2049809346;
assign addr[50945]= -2025707632;
assign addr[50946]= -1999036154;
assign addr[50947]= -1969828744;
assign addr[50948]= -1938122457;
assign addr[50949]= -1903957513;
assign addr[50950]= -1867377253;
assign addr[50951]= -1828428082;
assign addr[50952]= -1787159411;
assign addr[50953]= -1743623590;
assign addr[50954]= -1697875851;
assign addr[50955]= -1649974225;
assign addr[50956]= -1599979481;
assign addr[50957]= -1547955041;
assign addr[50958]= -1493966902;
assign addr[50959]= -1438083551;
assign addr[50960]= -1380375881;
assign addr[50961]= -1320917099;
assign addr[50962]= -1259782632;
assign addr[50963]= -1197050035;
assign addr[50964]= -1132798888;
assign addr[50965]= -1067110699;
assign addr[50966]= -1000068799;
assign addr[50967]= -931758235;
assign addr[50968]= -862265664;
assign addr[50969]= -791679244;
assign addr[50970]= -720088517;
assign addr[50971]= -647584304;
assign addr[50972]= -574258580;
assign addr[50973]= -500204365;
assign addr[50974]= -425515602;
assign addr[50975]= -350287041;
assign addr[50976]= -274614114;
assign addr[50977]= -198592817;
assign addr[50978]= -122319591;
assign addr[50979]= -45891193;
assign addr[50980]= 30595422;
assign addr[50981]= 107043224;
assign addr[50982]= 183355234;
assign addr[50983]= 259434643;
assign addr[50984]= 335184940;
assign addr[50985]= 410510029;
assign addr[50986]= 485314355;
assign addr[50987]= 559503022;
assign addr[50988]= 632981917;
assign addr[50989]= 705657826;
assign addr[50990]= 777438554;
assign addr[50991]= 848233042;
assign addr[50992]= 917951481;
assign addr[50993]= 986505429;
assign addr[50994]= 1053807919;
assign addr[50995]= 1119773573;
assign addr[50996]= 1184318708;
assign addr[50997]= 1247361445;
assign addr[50998]= 1308821808;
assign addr[50999]= 1368621831;
assign addr[51000]= 1426685652;
assign addr[51001]= 1482939614;
assign addr[51002]= 1537312353;
assign addr[51003]= 1589734894;
assign addr[51004]= 1640140734;
assign addr[51005]= 1688465931;
assign addr[51006]= 1734649179;
assign addr[51007]= 1778631892;
assign addr[51008]= 1820358275;
assign addr[51009]= 1859775393;
assign addr[51010]= 1896833245;
assign addr[51011]= 1931484818;
assign addr[51012]= 1963686155;
assign addr[51013]= 1993396407;
assign addr[51014]= 2020577882;
assign addr[51015]= 2045196100;
assign addr[51016]= 2067219829;
assign addr[51017]= 2086621133;
assign addr[51018]= 2103375398;
assign addr[51019]= 2117461370;
assign addr[51020]= 2128861181;
assign addr[51021]= 2137560369;
assign addr[51022]= 2143547897;
assign addr[51023]= 2146816171;
assign addr[51024]= 2147361045;
assign addr[51025]= 2145181827;
assign addr[51026]= 2140281282;
assign addr[51027]= 2132665626;
assign addr[51028]= 2122344521;
assign addr[51029]= 2109331059;
assign addr[51030]= 2093641749;
assign addr[51031]= 2075296495;
assign addr[51032]= 2054318569;
assign addr[51033]= 2030734582;
assign addr[51034]= 2004574453;
assign addr[51035]= 1975871368;
assign addr[51036]= 1944661739;
assign addr[51037]= 1910985158;
assign addr[51038]= 1874884346;
assign addr[51039]= 1836405100;
assign addr[51040]= 1795596234;
assign addr[51041]= 1752509516;
assign addr[51042]= 1707199606;
assign addr[51043]= 1659723983;
assign addr[51044]= 1610142873;
assign addr[51045]= 1558519173;
assign addr[51046]= 1504918373;
assign addr[51047]= 1449408469;
assign addr[51048]= 1392059879;
assign addr[51049]= 1332945355;
assign addr[51050]= 1272139887;
assign addr[51051]= 1209720613;
assign addr[51052]= 1145766716;
assign addr[51053]= 1080359326;
assign addr[51054]= 1013581418;
assign addr[51055]= 945517704;
assign addr[51056]= 876254528;
assign addr[51057]= 805879757;
assign addr[51058]= 734482665;
assign addr[51059]= 662153826;
assign addr[51060]= 588984994;
assign addr[51061]= 515068990;
assign addr[51062]= 440499581;
assign addr[51063]= 365371365;
assign addr[51064]= 289779648;
assign addr[51065]= 213820322;
assign addr[51066]= 137589750;
assign addr[51067]= 61184634;
assign addr[51068]= -15298099;
assign addr[51069]= -91761426;
assign addr[51070]= -168108346;
assign addr[51071]= -244242007;
assign addr[51072]= -320065829;
assign addr[51073]= -395483624;
assign addr[51074]= -470399716;
assign addr[51075]= -544719071;
assign addr[51076]= -618347408;
assign addr[51077]= -691191324;
assign addr[51078]= -763158411;
assign addr[51079]= -834157373;
assign addr[51080]= -904098143;
assign addr[51081]= -972891995;
assign addr[51082]= -1040451659;
assign addr[51083]= -1106691431;
assign addr[51084]= -1171527280;
assign addr[51085]= -1234876957;
assign addr[51086]= -1296660098;
assign addr[51087]= -1356798326;
assign addr[51088]= -1415215352;
assign addr[51089]= -1471837070;
assign addr[51090]= -1526591649;
assign addr[51091]= -1579409630;
assign addr[51092]= -1630224009;
assign addr[51093]= -1678970324;
assign addr[51094]= -1725586737;
assign addr[51095]= -1770014111;
assign addr[51096]= -1812196087;
assign addr[51097]= -1852079154;
assign addr[51098]= -1889612716;
assign addr[51099]= -1924749160;
assign addr[51100]= -1957443913;
assign addr[51101]= -1987655498;
assign addr[51102]= -2015345591;
assign addr[51103]= -2040479063;
assign addr[51104]= -2063024031;
assign addr[51105]= -2082951896;
assign addr[51106]= -2100237377;
assign addr[51107]= -2114858546;
assign addr[51108]= -2126796855;
assign addr[51109]= -2136037160;
assign addr[51110]= -2142567738;
assign addr[51111]= -2146380306;
assign addr[51112]= -2147470025;
assign addr[51113]= -2145835515;
assign addr[51114]= -2141478848;
assign addr[51115]= -2134405552;
assign addr[51116]= -2124624598;
assign addr[51117]= -2112148396;
assign addr[51118]= -2096992772;
assign addr[51119]= -2079176953;
assign addr[51120]= -2058723538;
assign addr[51121]= -2035658475;
assign addr[51122]= -2010011024;
assign addr[51123]= -1981813720;
assign addr[51124]= -1951102334;
assign addr[51125]= -1917915825;
assign addr[51126]= -1882296293;
assign addr[51127]= -1844288924;
assign addr[51128]= -1803941934;
assign addr[51129]= -1761306505;
assign addr[51130]= -1716436725;
assign addr[51131]= -1669389513;
assign addr[51132]= -1620224553;
assign addr[51133]= -1569004214;
assign addr[51134]= -1515793473;
assign addr[51135]= -1460659832;
assign addr[51136]= -1403673233;
assign addr[51137]= -1344905966;
assign addr[51138]= -1284432584;
assign addr[51139]= -1222329801;
assign addr[51140]= -1158676398;
assign addr[51141]= -1093553126;
assign addr[51142]= -1027042599;
assign addr[51143]= -959229189;
assign addr[51144]= -890198924;
assign addr[51145]= -820039373;
assign addr[51146]= -748839539;
assign addr[51147]= -676689746;
assign addr[51148]= -603681519;
assign addr[51149]= -529907477;
assign addr[51150]= -455461206;
assign addr[51151]= -380437148;
assign addr[51152]= -304930476;
assign addr[51153]= -229036977;
assign addr[51154]= -152852926;
assign addr[51155]= -76474970;
assign addr[51156]= 0;
assign addr[51157]= 76474970;
assign addr[51158]= 152852926;
assign addr[51159]= 229036977;
assign addr[51160]= 304930476;
assign addr[51161]= 380437148;
assign addr[51162]= 455461206;
assign addr[51163]= 529907477;
assign addr[51164]= 603681519;
assign addr[51165]= 676689746;
assign addr[51166]= 748839539;
assign addr[51167]= 820039373;
assign addr[51168]= 890198924;
assign addr[51169]= 959229189;
assign addr[51170]= 1027042599;
assign addr[51171]= 1093553126;
assign addr[51172]= 1158676398;
assign addr[51173]= 1222329801;
assign addr[51174]= 1284432584;
assign addr[51175]= 1344905966;
assign addr[51176]= 1403673233;
assign addr[51177]= 1460659832;
assign addr[51178]= 1515793473;
assign addr[51179]= 1569004214;
assign addr[51180]= 1620224553;
assign addr[51181]= 1669389513;
assign addr[51182]= 1716436725;
assign addr[51183]= 1761306505;
assign addr[51184]= 1803941934;
assign addr[51185]= 1844288924;
assign addr[51186]= 1882296293;
assign addr[51187]= 1917915825;
assign addr[51188]= 1951102334;
assign addr[51189]= 1981813720;
assign addr[51190]= 2010011024;
assign addr[51191]= 2035658475;
assign addr[51192]= 2058723538;
assign addr[51193]= 2079176953;
assign addr[51194]= 2096992772;
assign addr[51195]= 2112148396;
assign addr[51196]= 2124624598;
assign addr[51197]= 2134405552;
assign addr[51198]= 2141478848;
assign addr[51199]= 2145835515;
assign addr[51200]= 2147470025;
assign addr[51201]= 2146380306;
assign addr[51202]= 2142567738;
assign addr[51203]= 2136037160;
assign addr[51204]= 2126796855;
assign addr[51205]= 2114858546;
assign addr[51206]= 2100237377;
assign addr[51207]= 2082951896;
assign addr[51208]= 2063024031;
assign addr[51209]= 2040479063;
assign addr[51210]= 2015345591;
assign addr[51211]= 1987655498;
assign addr[51212]= 1957443913;
assign addr[51213]= 1924749160;
assign addr[51214]= 1889612716;
assign addr[51215]= 1852079154;
assign addr[51216]= 1812196087;
assign addr[51217]= 1770014111;
assign addr[51218]= 1725586737;
assign addr[51219]= 1678970324;
assign addr[51220]= 1630224009;
assign addr[51221]= 1579409630;
assign addr[51222]= 1526591649;
assign addr[51223]= 1471837070;
assign addr[51224]= 1415215352;
assign addr[51225]= 1356798326;
assign addr[51226]= 1296660098;
assign addr[51227]= 1234876957;
assign addr[51228]= 1171527280;
assign addr[51229]= 1106691431;
assign addr[51230]= 1040451659;
assign addr[51231]= 972891995;
assign addr[51232]= 904098143;
assign addr[51233]= 834157373;
assign addr[51234]= 763158411;
assign addr[51235]= 691191324;
assign addr[51236]= 618347408;
assign addr[51237]= 544719071;
assign addr[51238]= 470399716;
assign addr[51239]= 395483624;
assign addr[51240]= 320065829;
assign addr[51241]= 244242007;
assign addr[51242]= 168108346;
assign addr[51243]= 91761426;
assign addr[51244]= 15298099;
assign addr[51245]= -61184634;
assign addr[51246]= -137589750;
assign addr[51247]= -213820322;
assign addr[51248]= -289779648;
assign addr[51249]= -365371365;
assign addr[51250]= -440499581;
assign addr[51251]= -515068990;
assign addr[51252]= -588984994;
assign addr[51253]= -662153826;
assign addr[51254]= -734482665;
assign addr[51255]= -805879757;
assign addr[51256]= -876254528;
assign addr[51257]= -945517704;
assign addr[51258]= -1013581418;
assign addr[51259]= -1080359326;
assign addr[51260]= -1145766716;
assign addr[51261]= -1209720613;
assign addr[51262]= -1272139887;
assign addr[51263]= -1332945355;
assign addr[51264]= -1392059879;
assign addr[51265]= -1449408469;
assign addr[51266]= -1504918373;
assign addr[51267]= -1558519173;
assign addr[51268]= -1610142873;
assign addr[51269]= -1659723983;
assign addr[51270]= -1707199606;
assign addr[51271]= -1752509516;
assign addr[51272]= -1795596234;
assign addr[51273]= -1836405100;
assign addr[51274]= -1874884346;
assign addr[51275]= -1910985158;
assign addr[51276]= -1944661739;
assign addr[51277]= -1975871368;
assign addr[51278]= -2004574453;
assign addr[51279]= -2030734582;
assign addr[51280]= -2054318569;
assign addr[51281]= -2075296495;
assign addr[51282]= -2093641749;
assign addr[51283]= -2109331059;
assign addr[51284]= -2122344521;
assign addr[51285]= -2132665626;
assign addr[51286]= -2140281282;
assign addr[51287]= -2145181827;
assign addr[51288]= -2147361045;
assign addr[51289]= -2146816171;
assign addr[51290]= -2143547897;
assign addr[51291]= -2137560369;
assign addr[51292]= -2128861181;
assign addr[51293]= -2117461370;
assign addr[51294]= -2103375398;
assign addr[51295]= -2086621133;
assign addr[51296]= -2067219829;
assign addr[51297]= -2045196100;
assign addr[51298]= -2020577882;
assign addr[51299]= -1993396407;
assign addr[51300]= -1963686155;
assign addr[51301]= -1931484818;
assign addr[51302]= -1896833245;
assign addr[51303]= -1859775393;
assign addr[51304]= -1820358275;
assign addr[51305]= -1778631892;
assign addr[51306]= -1734649179;
assign addr[51307]= -1688465931;
assign addr[51308]= -1640140734;
assign addr[51309]= -1589734894;
assign addr[51310]= -1537312353;
assign addr[51311]= -1482939614;
assign addr[51312]= -1426685652;
assign addr[51313]= -1368621831;
assign addr[51314]= -1308821808;
assign addr[51315]= -1247361445;
assign addr[51316]= -1184318708;
assign addr[51317]= -1119773573;
assign addr[51318]= -1053807919;
assign addr[51319]= -986505429;
assign addr[51320]= -917951481;
assign addr[51321]= -848233042;
assign addr[51322]= -777438554;
assign addr[51323]= -705657826;
assign addr[51324]= -632981917;
assign addr[51325]= -559503022;
assign addr[51326]= -485314355;
assign addr[51327]= -410510029;
assign addr[51328]= -335184940;
assign addr[51329]= -259434643;
assign addr[51330]= -183355234;
assign addr[51331]= -107043224;
assign addr[51332]= -30595422;
assign addr[51333]= 45891193;
assign addr[51334]= 122319591;
assign addr[51335]= 198592817;
assign addr[51336]= 274614114;
assign addr[51337]= 350287041;
assign addr[51338]= 425515602;
assign addr[51339]= 500204365;
assign addr[51340]= 574258580;
assign addr[51341]= 647584304;
assign addr[51342]= 720088517;
assign addr[51343]= 791679244;
assign addr[51344]= 862265664;
assign addr[51345]= 931758235;
assign addr[51346]= 1000068799;
assign addr[51347]= 1067110699;
assign addr[51348]= 1132798888;
assign addr[51349]= 1197050035;
assign addr[51350]= 1259782632;
assign addr[51351]= 1320917099;
assign addr[51352]= 1380375881;
assign addr[51353]= 1438083551;
assign addr[51354]= 1493966902;
assign addr[51355]= 1547955041;
assign addr[51356]= 1599979481;
assign addr[51357]= 1649974225;
assign addr[51358]= 1697875851;
assign addr[51359]= 1743623590;
assign addr[51360]= 1787159411;
assign addr[51361]= 1828428082;
assign addr[51362]= 1867377253;
assign addr[51363]= 1903957513;
assign addr[51364]= 1938122457;
assign addr[51365]= 1969828744;
assign addr[51366]= 1999036154;
assign addr[51367]= 2025707632;
assign addr[51368]= 2049809346;
assign addr[51369]= 2071310720;
assign addr[51370]= 2090184478;
assign addr[51371]= 2106406677;
assign addr[51372]= 2119956737;
assign addr[51373]= 2130817471;
assign addr[51374]= 2138975100;
assign addr[51375]= 2144419275;
assign addr[51376]= 2147143090;
assign addr[51377]= 2147143090;
assign addr[51378]= 2144419275;
assign addr[51379]= 2138975100;
assign addr[51380]= 2130817471;
assign addr[51381]= 2119956737;
assign addr[51382]= 2106406677;
assign addr[51383]= 2090184478;
assign addr[51384]= 2071310720;
assign addr[51385]= 2049809346;
assign addr[51386]= 2025707632;
assign addr[51387]= 1999036154;
assign addr[51388]= 1969828744;
assign addr[51389]= 1938122457;
assign addr[51390]= 1903957513;
assign addr[51391]= 1867377253;
assign addr[51392]= 1828428082;
assign addr[51393]= 1787159411;
assign addr[51394]= 1743623590;
assign addr[51395]= 1697875851;
assign addr[51396]= 1649974225;
assign addr[51397]= 1599979481;
assign addr[51398]= 1547955041;
assign addr[51399]= 1493966902;
assign addr[51400]= 1438083551;
assign addr[51401]= 1380375881;
assign addr[51402]= 1320917099;
assign addr[51403]= 1259782632;
assign addr[51404]= 1197050035;
assign addr[51405]= 1132798888;
assign addr[51406]= 1067110699;
assign addr[51407]= 1000068799;
assign addr[51408]= 931758235;
assign addr[51409]= 862265664;
assign addr[51410]= 791679244;
assign addr[51411]= 720088517;
assign addr[51412]= 647584304;
assign addr[51413]= 574258580;
assign addr[51414]= 500204365;
assign addr[51415]= 425515602;
assign addr[51416]= 350287041;
assign addr[51417]= 274614114;
assign addr[51418]= 198592817;
assign addr[51419]= 122319591;
assign addr[51420]= 45891193;
assign addr[51421]= -30595422;
assign addr[51422]= -107043224;
assign addr[51423]= -183355234;
assign addr[51424]= -259434643;
assign addr[51425]= -335184940;
assign addr[51426]= -410510029;
assign addr[51427]= -485314355;
assign addr[51428]= -559503022;
assign addr[51429]= -632981917;
assign addr[51430]= -705657826;
assign addr[51431]= -777438554;
assign addr[51432]= -848233042;
assign addr[51433]= -917951481;
assign addr[51434]= -986505429;
assign addr[51435]= -1053807919;
assign addr[51436]= -1119773573;
assign addr[51437]= -1184318708;
assign addr[51438]= -1247361445;
assign addr[51439]= -1308821808;
assign addr[51440]= -1368621831;
assign addr[51441]= -1426685652;
assign addr[51442]= -1482939614;
assign addr[51443]= -1537312353;
assign addr[51444]= -1589734894;
assign addr[51445]= -1640140734;
assign addr[51446]= -1688465931;
assign addr[51447]= -1734649179;
assign addr[51448]= -1778631892;
assign addr[51449]= -1820358275;
assign addr[51450]= -1859775393;
assign addr[51451]= -1896833245;
assign addr[51452]= -1931484818;
assign addr[51453]= -1963686155;
assign addr[51454]= -1993396407;
assign addr[51455]= -2020577882;
assign addr[51456]= -2045196100;
assign addr[51457]= -2067219829;
assign addr[51458]= -2086621133;
assign addr[51459]= -2103375398;
assign addr[51460]= -2117461370;
assign addr[51461]= -2128861181;
assign addr[51462]= -2137560369;
assign addr[51463]= -2143547897;
assign addr[51464]= -2146816171;
assign addr[51465]= -2147361045;
assign addr[51466]= -2145181827;
assign addr[51467]= -2140281282;
assign addr[51468]= -2132665626;
assign addr[51469]= -2122344521;
assign addr[51470]= -2109331059;
assign addr[51471]= -2093641749;
assign addr[51472]= -2075296495;
assign addr[51473]= -2054318569;
assign addr[51474]= -2030734582;
assign addr[51475]= -2004574453;
assign addr[51476]= -1975871368;
assign addr[51477]= -1944661739;
assign addr[51478]= -1910985158;
assign addr[51479]= -1874884346;
assign addr[51480]= -1836405100;
assign addr[51481]= -1795596234;
assign addr[51482]= -1752509516;
assign addr[51483]= -1707199606;
assign addr[51484]= -1659723983;
assign addr[51485]= -1610142873;
assign addr[51486]= -1558519173;
assign addr[51487]= -1504918373;
assign addr[51488]= -1449408469;
assign addr[51489]= -1392059879;
assign addr[51490]= -1332945355;
assign addr[51491]= -1272139887;
assign addr[51492]= -1209720613;
assign addr[51493]= -1145766716;
assign addr[51494]= -1080359326;
assign addr[51495]= -1013581418;
assign addr[51496]= -945517704;
assign addr[51497]= -876254528;
assign addr[51498]= -805879757;
assign addr[51499]= -734482665;
assign addr[51500]= -662153826;
assign addr[51501]= -588984994;
assign addr[51502]= -515068990;
assign addr[51503]= -440499581;
assign addr[51504]= -365371365;
assign addr[51505]= -289779648;
assign addr[51506]= -213820322;
assign addr[51507]= -137589750;
assign addr[51508]= -61184634;
assign addr[51509]= 15298099;
assign addr[51510]= 91761426;
assign addr[51511]= 168108346;
assign addr[51512]= 244242007;
assign addr[51513]= 320065829;
assign addr[51514]= 395483624;
assign addr[51515]= 470399716;
assign addr[51516]= 544719071;
assign addr[51517]= 618347408;
assign addr[51518]= 691191324;
assign addr[51519]= 763158411;
assign addr[51520]= 834157373;
assign addr[51521]= 904098143;
assign addr[51522]= 972891995;
assign addr[51523]= 1040451659;
assign addr[51524]= 1106691431;
assign addr[51525]= 1171527280;
assign addr[51526]= 1234876957;
assign addr[51527]= 1296660098;
assign addr[51528]= 1356798326;
assign addr[51529]= 1415215352;
assign addr[51530]= 1471837070;
assign addr[51531]= 1526591649;
assign addr[51532]= 1579409630;
assign addr[51533]= 1630224009;
assign addr[51534]= 1678970324;
assign addr[51535]= 1725586737;
assign addr[51536]= 1770014111;
assign addr[51537]= 1812196087;
assign addr[51538]= 1852079154;
assign addr[51539]= 1889612716;
assign addr[51540]= 1924749160;
assign addr[51541]= 1957443913;
assign addr[51542]= 1987655498;
assign addr[51543]= 2015345591;
assign addr[51544]= 2040479063;
assign addr[51545]= 2063024031;
assign addr[51546]= 2082951896;
assign addr[51547]= 2100237377;
assign addr[51548]= 2114858546;
assign addr[51549]= 2126796855;
assign addr[51550]= 2136037160;
assign addr[51551]= 2142567738;
assign addr[51552]= 2146380306;
assign addr[51553]= 2147470025;
assign addr[51554]= 2145835515;
assign addr[51555]= 2141478848;
assign addr[51556]= 2134405552;
assign addr[51557]= 2124624598;
assign addr[51558]= 2112148396;
assign addr[51559]= 2096992772;
assign addr[51560]= 2079176953;
assign addr[51561]= 2058723538;
assign addr[51562]= 2035658475;
assign addr[51563]= 2010011024;
assign addr[51564]= 1981813720;
assign addr[51565]= 1951102334;
assign addr[51566]= 1917915825;
assign addr[51567]= 1882296293;
assign addr[51568]= 1844288924;
assign addr[51569]= 1803941934;
assign addr[51570]= 1761306505;
assign addr[51571]= 1716436725;
assign addr[51572]= 1669389513;
assign addr[51573]= 1620224553;
assign addr[51574]= 1569004214;
assign addr[51575]= 1515793473;
assign addr[51576]= 1460659832;
assign addr[51577]= 1403673233;
assign addr[51578]= 1344905966;
assign addr[51579]= 1284432584;
assign addr[51580]= 1222329801;
assign addr[51581]= 1158676398;
assign addr[51582]= 1093553126;
assign addr[51583]= 1027042599;
assign addr[51584]= 959229189;
assign addr[51585]= 890198924;
assign addr[51586]= 820039373;
assign addr[51587]= 748839539;
assign addr[51588]= 676689746;
assign addr[51589]= 603681519;
assign addr[51590]= 529907477;
assign addr[51591]= 455461206;
assign addr[51592]= 380437148;
assign addr[51593]= 304930476;
assign addr[51594]= 229036977;
assign addr[51595]= 152852926;
assign addr[51596]= 76474970;
assign addr[51597]= 0;
assign addr[51598]= -76474970;
assign addr[51599]= -152852926;
assign addr[51600]= -229036977;
assign addr[51601]= -304930476;
assign addr[51602]= -380437148;
assign addr[51603]= -455461206;
assign addr[51604]= -529907477;
assign addr[51605]= -603681519;
assign addr[51606]= -676689746;
assign addr[51607]= -748839539;
assign addr[51608]= -820039373;
assign addr[51609]= -890198924;
assign addr[51610]= -959229189;
assign addr[51611]= -1027042599;
assign addr[51612]= -1093553126;
assign addr[51613]= -1158676398;
assign addr[51614]= -1222329801;
assign addr[51615]= -1284432584;
assign addr[51616]= -1344905966;
assign addr[51617]= -1403673233;
assign addr[51618]= -1460659832;
assign addr[51619]= -1515793473;
assign addr[51620]= -1569004214;
assign addr[51621]= -1620224553;
assign addr[51622]= -1669389513;
assign addr[51623]= -1716436725;
assign addr[51624]= -1761306505;
assign addr[51625]= -1803941934;
assign addr[51626]= -1844288924;
assign addr[51627]= -1882296293;
assign addr[51628]= -1917915825;
assign addr[51629]= -1951102334;
assign addr[51630]= -1981813720;
assign addr[51631]= -2010011024;
assign addr[51632]= -2035658475;
assign addr[51633]= -2058723538;
assign addr[51634]= -2079176953;
assign addr[51635]= -2096992772;
assign addr[51636]= -2112148396;
assign addr[51637]= -2124624598;
assign addr[51638]= -2134405552;
assign addr[51639]= -2141478848;
assign addr[51640]= -2145835515;
assign addr[51641]= -2147470025;
assign addr[51642]= -2146380306;
assign addr[51643]= -2142567738;
assign addr[51644]= -2136037160;
assign addr[51645]= -2126796855;
assign addr[51646]= -2114858546;
assign addr[51647]= -2100237377;
assign addr[51648]= -2082951896;
assign addr[51649]= -2063024031;
assign addr[51650]= -2040479063;
assign addr[51651]= -2015345591;
assign addr[51652]= -1987655498;
assign addr[51653]= -1957443913;
assign addr[51654]= -1924749160;
assign addr[51655]= -1889612716;
assign addr[51656]= -1852079154;
assign addr[51657]= -1812196087;
assign addr[51658]= -1770014111;
assign addr[51659]= -1725586737;
assign addr[51660]= -1678970324;
assign addr[51661]= -1630224009;
assign addr[51662]= -1579409630;
assign addr[51663]= -1526591649;
assign addr[51664]= -1471837070;
assign addr[51665]= -1415215352;
assign addr[51666]= -1356798326;
assign addr[51667]= -1296660098;
assign addr[51668]= -1234876957;
assign addr[51669]= -1171527280;
assign addr[51670]= -1106691431;
assign addr[51671]= -1040451659;
assign addr[51672]= -972891995;
assign addr[51673]= -904098143;
assign addr[51674]= -834157373;
assign addr[51675]= -763158411;
assign addr[51676]= -691191324;
assign addr[51677]= -618347408;
assign addr[51678]= -544719071;
assign addr[51679]= -470399716;
assign addr[51680]= -395483624;
assign addr[51681]= -320065829;
assign addr[51682]= -244242007;
assign addr[51683]= -168108346;
assign addr[51684]= -91761426;
assign addr[51685]= -15298099;
assign addr[51686]= 61184634;
assign addr[51687]= 137589750;
assign addr[51688]= 213820322;
assign addr[51689]= 289779648;
assign addr[51690]= 365371365;
assign addr[51691]= 440499581;
assign addr[51692]= 515068990;
assign addr[51693]= 588984994;
assign addr[51694]= 662153826;
assign addr[51695]= 734482665;
assign addr[51696]= 805879757;
assign addr[51697]= 876254528;
assign addr[51698]= 945517704;
assign addr[51699]= 1013581418;
assign addr[51700]= 1080359326;
assign addr[51701]= 1145766716;
assign addr[51702]= 1209720613;
assign addr[51703]= 1272139887;
assign addr[51704]= 1332945355;
assign addr[51705]= 1392059879;
assign addr[51706]= 1449408469;
assign addr[51707]= 1504918373;
assign addr[51708]= 1558519173;
assign addr[51709]= 1610142873;
assign addr[51710]= 1659723983;
assign addr[51711]= 1707199606;
assign addr[51712]= 1752509516;
assign addr[51713]= 1795596234;
assign addr[51714]= 1836405100;
assign addr[51715]= 1874884346;
assign addr[51716]= 1910985158;
assign addr[51717]= 1944661739;
assign addr[51718]= 1975871368;
assign addr[51719]= 2004574453;
assign addr[51720]= 2030734582;
assign addr[51721]= 2054318569;
assign addr[51722]= 2075296495;
assign addr[51723]= 2093641749;
assign addr[51724]= 2109331059;
assign addr[51725]= 2122344521;
assign addr[51726]= 2132665626;
assign addr[51727]= 2140281282;
assign addr[51728]= 2145181827;
assign addr[51729]= 2147361045;
assign addr[51730]= 2146816171;
assign addr[51731]= 2143547897;
assign addr[51732]= 2137560369;
assign addr[51733]= 2128861181;
assign addr[51734]= 2117461370;
assign addr[51735]= 2103375398;
assign addr[51736]= 2086621133;
assign addr[51737]= 2067219829;
assign addr[51738]= 2045196100;
assign addr[51739]= 2020577882;
assign addr[51740]= 1993396407;
assign addr[51741]= 1963686155;
assign addr[51742]= 1931484818;
assign addr[51743]= 1896833245;
assign addr[51744]= 1859775393;
assign addr[51745]= 1820358275;
assign addr[51746]= 1778631892;
assign addr[51747]= 1734649179;
assign addr[51748]= 1688465931;
assign addr[51749]= 1640140734;
assign addr[51750]= 1589734894;
assign addr[51751]= 1537312353;
assign addr[51752]= 1482939614;
assign addr[51753]= 1426685652;
assign addr[51754]= 1368621831;
assign addr[51755]= 1308821808;
assign addr[51756]= 1247361445;
assign addr[51757]= 1184318708;
assign addr[51758]= 1119773573;
assign addr[51759]= 1053807919;
assign addr[51760]= 986505429;
assign addr[51761]= 917951481;
assign addr[51762]= 848233042;
assign addr[51763]= 777438554;
assign addr[51764]= 705657826;
assign addr[51765]= 632981917;
assign addr[51766]= 559503022;
assign addr[51767]= 485314355;
assign addr[51768]= 410510029;
assign addr[51769]= 335184940;
assign addr[51770]= 259434643;
assign addr[51771]= 183355234;
assign addr[51772]= 107043224;
assign addr[51773]= 30595422;
assign addr[51774]= -45891193;
assign addr[51775]= -122319591;
assign addr[51776]= -198592817;
assign addr[51777]= -274614114;
assign addr[51778]= -350287041;
assign addr[51779]= -425515602;
assign addr[51780]= -500204365;
assign addr[51781]= -574258580;
assign addr[51782]= -647584304;
assign addr[51783]= -720088517;
assign addr[51784]= -791679244;
assign addr[51785]= -862265664;
assign addr[51786]= -931758235;
assign addr[51787]= -1000068799;
assign addr[51788]= -1067110699;
assign addr[51789]= -1132798888;
assign addr[51790]= -1197050035;
assign addr[51791]= -1259782632;
assign addr[51792]= -1320917099;
assign addr[51793]= -1380375881;
assign addr[51794]= -1438083551;
assign addr[51795]= -1493966902;
assign addr[51796]= -1547955041;
assign addr[51797]= -1599979481;
assign addr[51798]= -1649974225;
assign addr[51799]= -1697875851;
assign addr[51800]= -1743623590;
assign addr[51801]= -1787159411;
assign addr[51802]= -1828428082;
assign addr[51803]= -1867377253;
assign addr[51804]= -1903957513;
assign addr[51805]= -1938122457;
assign addr[51806]= -1969828744;
assign addr[51807]= -1999036154;
assign addr[51808]= -2025707632;
assign addr[51809]= -2049809346;
assign addr[51810]= -2071310720;
assign addr[51811]= -2090184478;
assign addr[51812]= -2106406677;
assign addr[51813]= -2119956737;
assign addr[51814]= -2130817471;
assign addr[51815]= -2138975100;
assign addr[51816]= -2144419275;
assign addr[51817]= -2147143090;
assign addr[51818]= -2147143090;
assign addr[51819]= -2144419275;
assign addr[51820]= -2138975100;
assign addr[51821]= -2130817471;
assign addr[51822]= -2119956737;
assign addr[51823]= -2106406677;
assign addr[51824]= -2090184478;
assign addr[51825]= -2071310720;
assign addr[51826]= -2049809346;
assign addr[51827]= -2025707632;
assign addr[51828]= -1999036154;
assign addr[51829]= -1969828744;
assign addr[51830]= -1938122457;
assign addr[51831]= -1903957513;
assign addr[51832]= -1867377253;
assign addr[51833]= -1828428082;
assign addr[51834]= -1787159411;
assign addr[51835]= -1743623590;
assign addr[51836]= -1697875851;
assign addr[51837]= -1649974225;
assign addr[51838]= -1599979481;
assign addr[51839]= -1547955041;
assign addr[51840]= -1493966902;
assign addr[51841]= -1438083551;
assign addr[51842]= -1380375881;
assign addr[51843]= -1320917099;
assign addr[51844]= -1259782632;
assign addr[51845]= -1197050035;
assign addr[51846]= -1132798888;
assign addr[51847]= -1067110699;
assign addr[51848]= -1000068799;
assign addr[51849]= -931758235;
assign addr[51850]= -862265664;
assign addr[51851]= -791679244;
assign addr[51852]= -720088517;
assign addr[51853]= -647584304;
assign addr[51854]= -574258580;
assign addr[51855]= -500204365;
assign addr[51856]= -425515602;
assign addr[51857]= -350287041;
assign addr[51858]= -274614114;
assign addr[51859]= -198592817;
assign addr[51860]= -122319591;
assign addr[51861]= -45891193;
assign addr[51862]= 30595422;
assign addr[51863]= 107043224;
assign addr[51864]= 183355234;
assign addr[51865]= 259434643;
assign addr[51866]= 335184940;
assign addr[51867]= 410510029;
assign addr[51868]= 485314355;
assign addr[51869]= 559503022;
assign addr[51870]= 632981917;
assign addr[51871]= 705657826;
assign addr[51872]= 777438554;
assign addr[51873]= 848233042;
assign addr[51874]= 917951481;
assign addr[51875]= 986505429;
assign addr[51876]= 1053807919;
assign addr[51877]= 1119773573;
assign addr[51878]= 1184318708;
assign addr[51879]= 1247361445;
assign addr[51880]= 1308821808;
assign addr[51881]= 1368621831;
assign addr[51882]= 1426685652;
assign addr[51883]= 1482939614;
assign addr[51884]= 1537312353;
assign addr[51885]= 1589734894;
assign addr[51886]= 1640140734;
assign addr[51887]= 1688465931;
assign addr[51888]= 1734649179;
assign addr[51889]= 1778631892;
assign addr[51890]= 1820358275;
assign addr[51891]= 1859775393;
assign addr[51892]= 1896833245;
assign addr[51893]= 1931484818;
assign addr[51894]= 1963686155;
assign addr[51895]= 1993396407;
assign addr[51896]= 2020577882;
assign addr[51897]= 2045196100;
assign addr[51898]= 2067219829;
assign addr[51899]= 2086621133;
assign addr[51900]= 2103375398;
assign addr[51901]= 2117461370;
assign addr[51902]= 2128861181;
assign addr[51903]= 2137560369;
assign addr[51904]= 2143547897;
assign addr[51905]= 2146816171;
assign addr[51906]= 2147361045;
assign addr[51907]= 2145181827;
assign addr[51908]= 2140281282;
assign addr[51909]= 2132665626;
assign addr[51910]= 2122344521;
assign addr[51911]= 2109331059;
assign addr[51912]= 2093641749;
assign addr[51913]= 2075296495;
assign addr[51914]= 2054318569;
assign addr[51915]= 2030734582;
assign addr[51916]= 2004574453;
assign addr[51917]= 1975871368;
assign addr[51918]= 1944661739;
assign addr[51919]= 1910985158;
assign addr[51920]= 1874884346;
assign addr[51921]= 1836405100;
assign addr[51922]= 1795596234;
assign addr[51923]= 1752509516;
assign addr[51924]= 1707199606;
assign addr[51925]= 1659723983;
assign addr[51926]= 1610142873;
assign addr[51927]= 1558519173;
assign addr[51928]= 1504918373;
assign addr[51929]= 1449408469;
assign addr[51930]= 1392059879;
assign addr[51931]= 1332945355;
assign addr[51932]= 1272139887;
assign addr[51933]= 1209720613;
assign addr[51934]= 1145766716;
assign addr[51935]= 1080359326;
assign addr[51936]= 1013581418;
assign addr[51937]= 945517704;
assign addr[51938]= 876254528;
assign addr[51939]= 805879757;
assign addr[51940]= 734482665;
assign addr[51941]= 662153826;
assign addr[51942]= 588984994;
assign addr[51943]= 515068990;
assign addr[51944]= 440499581;
assign addr[51945]= 365371365;
assign addr[51946]= 289779648;
assign addr[51947]= 213820322;
assign addr[51948]= 137589750;
assign addr[51949]= 61184634;
assign addr[51950]= -15298099;
assign addr[51951]= -91761426;
assign addr[51952]= -168108346;
assign addr[51953]= -244242007;
assign addr[51954]= -320065829;
assign addr[51955]= -395483624;
assign addr[51956]= -470399716;
assign addr[51957]= -544719071;
assign addr[51958]= -618347408;
assign addr[51959]= -691191324;
assign addr[51960]= -763158411;
assign addr[51961]= -834157373;
assign addr[51962]= -904098143;
assign addr[51963]= -972891995;
assign addr[51964]= -1040451659;
assign addr[51965]= -1106691431;
assign addr[51966]= -1171527280;
assign addr[51967]= -1234876957;
assign addr[51968]= -1296660098;
assign addr[51969]= -1356798326;
assign addr[51970]= -1415215352;
assign addr[51971]= -1471837070;
assign addr[51972]= -1526591649;
assign addr[51973]= -1579409630;
assign addr[51974]= -1630224009;
assign addr[51975]= -1678970324;
assign addr[51976]= -1725586737;
assign addr[51977]= -1770014111;
assign addr[51978]= -1812196087;
assign addr[51979]= -1852079154;
assign addr[51980]= -1889612716;
assign addr[51981]= -1924749160;
assign addr[51982]= -1957443913;
assign addr[51983]= -1987655498;
assign addr[51984]= -2015345591;
assign addr[51985]= -2040479063;
assign addr[51986]= -2063024031;
assign addr[51987]= -2082951896;
assign addr[51988]= -2100237377;
assign addr[51989]= -2114858546;
assign addr[51990]= -2126796855;
assign addr[51991]= -2136037160;
assign addr[51992]= -2142567738;
assign addr[51993]= -2146380306;
assign addr[51994]= -2147470025;
assign addr[51995]= -2145835515;
assign addr[51996]= -2141478848;
assign addr[51997]= -2134405552;
assign addr[51998]= -2124624598;
assign addr[51999]= -2112148396;
assign addr[52000]= -2096992772;
assign addr[52001]= -2079176953;
assign addr[52002]= -2058723538;
assign addr[52003]= -2035658475;
assign addr[52004]= -2010011024;
assign addr[52005]= -1981813720;
assign addr[52006]= -1951102334;
assign addr[52007]= -1917915825;
assign addr[52008]= -1882296293;
assign addr[52009]= -1844288924;
assign addr[52010]= -1803941934;
assign addr[52011]= -1761306505;
assign addr[52012]= -1716436725;
assign addr[52013]= -1669389513;
assign addr[52014]= -1620224553;
assign addr[52015]= -1569004214;
assign addr[52016]= -1515793473;
assign addr[52017]= -1460659832;
assign addr[52018]= -1403673233;
assign addr[52019]= -1344905966;
assign addr[52020]= -1284432584;
assign addr[52021]= -1222329801;
assign addr[52022]= -1158676398;
assign addr[52023]= -1093553126;
assign addr[52024]= -1027042599;
assign addr[52025]= -959229189;
assign addr[52026]= -890198924;
assign addr[52027]= -820039373;
assign addr[52028]= -748839539;
assign addr[52029]= -676689746;
assign addr[52030]= -603681519;
assign addr[52031]= -529907477;
assign addr[52032]= -455461206;
assign addr[52033]= -380437148;
assign addr[52034]= -304930476;
assign addr[52035]= -229036977;
assign addr[52036]= -152852926;
assign addr[52037]= -76474970;
assign addr[52038]= 0;
assign addr[52039]= 76474970;
assign addr[52040]= 152852926;
assign addr[52041]= 229036977;
assign addr[52042]= 304930476;
assign addr[52043]= 380437148;
assign addr[52044]= 455461206;
assign addr[52045]= 529907477;
assign addr[52046]= 603681519;
assign addr[52047]= 676689746;
assign addr[52048]= 748839539;
assign addr[52049]= 820039373;
assign addr[52050]= 890198924;
assign addr[52051]= 959229189;
assign addr[52052]= 1027042599;
assign addr[52053]= 1093553126;
assign addr[52054]= 1158676398;
assign addr[52055]= 1222329801;
assign addr[52056]= 1284432584;
assign addr[52057]= 1344905966;
assign addr[52058]= 1403673233;
assign addr[52059]= 1460659832;
assign addr[52060]= 1515793473;
assign addr[52061]= 1569004214;
assign addr[52062]= 1620224553;
assign addr[52063]= 1669389513;
assign addr[52064]= 1716436725;
assign addr[52065]= 1761306505;
assign addr[52066]= 1803941934;
assign addr[52067]= 1844288924;
assign addr[52068]= 1882296293;
assign addr[52069]= 1917915825;
assign addr[52070]= 1951102334;
assign addr[52071]= 1981813720;
assign addr[52072]= 2010011024;
assign addr[52073]= 2035658475;
assign addr[52074]= 2058723538;
assign addr[52075]= 2079176953;
assign addr[52076]= 2096992772;
assign addr[52077]= 2112148396;
assign addr[52078]= 2124624598;
assign addr[52079]= 2134405552;
assign addr[52080]= 2141478848;
assign addr[52081]= 2145835515;
assign addr[52082]= 2147470025;
assign addr[52083]= 2146380306;
assign addr[52084]= 2142567738;
assign addr[52085]= 2136037160;
assign addr[52086]= 2126796855;
assign addr[52087]= 2114858546;
assign addr[52088]= 2100237377;
assign addr[52089]= 2082951896;
assign addr[52090]= 2063024031;
assign addr[52091]= 2040479063;
assign addr[52092]= 2015345591;
assign addr[52093]= 1987655498;
assign addr[52094]= 1957443913;
assign addr[52095]= 1924749160;
assign addr[52096]= 1889612716;
assign addr[52097]= 1852079154;
assign addr[52098]= 1812196087;
assign addr[52099]= 1770014111;
assign addr[52100]= 1725586737;
assign addr[52101]= 1678970324;
assign addr[52102]= 1630224009;
assign addr[52103]= 1579409630;
assign addr[52104]= 1526591649;
assign addr[52105]= 1471837070;
assign addr[52106]= 1415215352;
assign addr[52107]= 1356798326;
assign addr[52108]= 1296660098;
assign addr[52109]= 1234876957;
assign addr[52110]= 1171527280;
assign addr[52111]= 1106691431;
assign addr[52112]= 1040451659;
assign addr[52113]= 972891995;
assign addr[52114]= 904098143;
assign addr[52115]= 834157373;
assign addr[52116]= 763158411;
assign addr[52117]= 691191324;
assign addr[52118]= 618347408;
assign addr[52119]= 544719071;
assign addr[52120]= 470399716;
assign addr[52121]= 395483624;
assign addr[52122]= 320065829;
assign addr[52123]= 244242007;
assign addr[52124]= 168108346;
assign addr[52125]= 91761426;
assign addr[52126]= 15298099;
assign addr[52127]= -61184634;
assign addr[52128]= -137589750;
assign addr[52129]= -213820322;
assign addr[52130]= -289779648;
assign addr[52131]= -365371365;
assign addr[52132]= -440499581;
assign addr[52133]= -515068990;
assign addr[52134]= -588984994;
assign addr[52135]= -662153826;
assign addr[52136]= -734482665;
assign addr[52137]= -805879757;
assign addr[52138]= -876254528;
assign addr[52139]= -945517704;
assign addr[52140]= -1013581418;
assign addr[52141]= -1080359326;
assign addr[52142]= -1145766716;
assign addr[52143]= -1209720613;
assign addr[52144]= -1272139887;
assign addr[52145]= -1332945355;
assign addr[52146]= -1392059879;
assign addr[52147]= -1449408469;
assign addr[52148]= -1504918373;
assign addr[52149]= -1558519173;
assign addr[52150]= -1610142873;
assign addr[52151]= -1659723983;
assign addr[52152]= -1707199606;
assign addr[52153]= -1752509516;
assign addr[52154]= -1795596234;
assign addr[52155]= -1836405100;
assign addr[52156]= -1874884346;
assign addr[52157]= -1910985158;
assign addr[52158]= -1944661739;
assign addr[52159]= -1975871368;
assign addr[52160]= -2004574453;
assign addr[52161]= -2030734582;
assign addr[52162]= -2054318569;
assign addr[52163]= -2075296495;
assign addr[52164]= -2093641749;
assign addr[52165]= -2109331059;
assign addr[52166]= -2122344521;
assign addr[52167]= -2132665626;
assign addr[52168]= -2140281282;
assign addr[52169]= -2145181827;
assign addr[52170]= -2147361045;
assign addr[52171]= -2146816171;
assign addr[52172]= -2143547897;
assign addr[52173]= -2137560369;
assign addr[52174]= -2128861181;
assign addr[52175]= -2117461370;
assign addr[52176]= -2103375398;
assign addr[52177]= -2086621133;
assign addr[52178]= -2067219829;
assign addr[52179]= -2045196100;
assign addr[52180]= -2020577882;
assign addr[52181]= -1993396407;
assign addr[52182]= -1963686155;
assign addr[52183]= -1931484818;
assign addr[52184]= -1896833245;
assign addr[52185]= -1859775393;
assign addr[52186]= -1820358275;
assign addr[52187]= -1778631892;
assign addr[52188]= -1734649179;
assign addr[52189]= -1688465931;
assign addr[52190]= -1640140734;
assign addr[52191]= -1589734894;
assign addr[52192]= -1537312353;
assign addr[52193]= -1482939614;
assign addr[52194]= -1426685652;
assign addr[52195]= -1368621831;
assign addr[52196]= -1308821808;
assign addr[52197]= -1247361445;
assign addr[52198]= -1184318708;
assign addr[52199]= -1119773573;
assign addr[52200]= -1053807919;
assign addr[52201]= -986505429;
assign addr[52202]= -917951481;
assign addr[52203]= -848233042;
assign addr[52204]= -777438554;
assign addr[52205]= -705657826;
assign addr[52206]= -632981917;
assign addr[52207]= -559503022;
assign addr[52208]= -485314355;
assign addr[52209]= -410510029;
assign addr[52210]= -335184940;
assign addr[52211]= -259434643;
assign addr[52212]= -183355234;
assign addr[52213]= -107043224;
assign addr[52214]= -30595422;
assign addr[52215]= 45891193;
assign addr[52216]= 122319591;
assign addr[52217]= 198592817;
assign addr[52218]= 274614114;
assign addr[52219]= 350287041;
assign addr[52220]= 425515602;
assign addr[52221]= 500204365;
assign addr[52222]= 574258580;
assign addr[52223]= 647584304;
assign addr[52224]= 720088517;
assign addr[52225]= 791679244;
assign addr[52226]= 862265664;
assign addr[52227]= 931758235;
assign addr[52228]= 1000068799;
assign addr[52229]= 1067110699;
assign addr[52230]= 1132798888;
assign addr[52231]= 1197050035;
assign addr[52232]= 1259782632;
assign addr[52233]= 1320917099;
assign addr[52234]= 1380375881;
assign addr[52235]= 1438083551;
assign addr[52236]= 1493966902;
assign addr[52237]= 1547955041;
assign addr[52238]= 1599979481;
assign addr[52239]= 1649974225;
assign addr[52240]= 1697875851;
assign addr[52241]= 1743623590;
assign addr[52242]= 1787159411;
assign addr[52243]= 1828428082;
assign addr[52244]= 1867377253;
assign addr[52245]= 1903957513;
assign addr[52246]= 1938122457;
assign addr[52247]= 1969828744;
assign addr[52248]= 1999036154;
assign addr[52249]= 2025707632;
assign addr[52250]= 2049809346;
assign addr[52251]= 2071310720;
assign addr[52252]= 2090184478;
assign addr[52253]= 2106406677;
assign addr[52254]= 2119956737;
assign addr[52255]= 2130817471;
assign addr[52256]= 2138975100;
assign addr[52257]= 2144419275;
assign addr[52258]= 2147143090;
assign addr[52259]= 2147143090;
assign addr[52260]= 2144419275;
assign addr[52261]= 2138975100;
assign addr[52262]= 2130817471;
assign addr[52263]= 2119956737;
assign addr[52264]= 2106406677;
assign addr[52265]= 2090184478;
assign addr[52266]= 2071310720;
assign addr[52267]= 2049809346;
assign addr[52268]= 2025707632;
assign addr[52269]= 1999036154;
assign addr[52270]= 1969828744;
assign addr[52271]= 1938122457;
assign addr[52272]= 1903957513;
assign addr[52273]= 1867377253;
assign addr[52274]= 1828428082;
assign addr[52275]= 1787159411;
assign addr[52276]= 1743623590;
assign addr[52277]= 1697875851;
assign addr[52278]= 1649974225;
assign addr[52279]= 1599979481;
assign addr[52280]= 1547955041;
assign addr[52281]= 1493966902;
assign addr[52282]= 1438083551;
assign addr[52283]= 1380375881;
assign addr[52284]= 1320917099;
assign addr[52285]= 1259782632;
assign addr[52286]= 1197050035;
assign addr[52287]= 1132798888;
assign addr[52288]= 1067110699;
assign addr[52289]= 1000068799;
assign addr[52290]= 931758235;
assign addr[52291]= 862265664;
assign addr[52292]= 791679244;
assign addr[52293]= 720088517;
assign addr[52294]= 647584304;
assign addr[52295]= 574258580;
assign addr[52296]= 500204365;
assign addr[52297]= 425515602;
assign addr[52298]= 350287041;
assign addr[52299]= 274614114;
assign addr[52300]= 198592817;
assign addr[52301]= 122319591;
assign addr[52302]= 45891193;
assign addr[52303]= -30595422;
assign addr[52304]= -107043224;
assign addr[52305]= -183355234;
assign addr[52306]= -259434643;
assign addr[52307]= -335184940;
assign addr[52308]= -410510029;
assign addr[52309]= -485314355;
assign addr[52310]= -559503022;
assign addr[52311]= -632981917;
assign addr[52312]= -705657826;
assign addr[52313]= -777438554;
assign addr[52314]= -848233042;
assign addr[52315]= -917951481;
assign addr[52316]= -986505429;
assign addr[52317]= -1053807919;
assign addr[52318]= -1119773573;
assign addr[52319]= -1184318708;
assign addr[52320]= -1247361445;
assign addr[52321]= -1308821808;
assign addr[52322]= -1368621831;
assign addr[52323]= -1426685652;
assign addr[52324]= -1482939614;
assign addr[52325]= -1537312353;
assign addr[52326]= -1589734894;
assign addr[52327]= -1640140734;
assign addr[52328]= -1688465931;
assign addr[52329]= -1734649179;
assign addr[52330]= -1778631892;
assign addr[52331]= -1820358275;
assign addr[52332]= -1859775393;
assign addr[52333]= -1896833245;
assign addr[52334]= -1931484818;
assign addr[52335]= -1963686155;
assign addr[52336]= -1993396407;
assign addr[52337]= -2020577882;
assign addr[52338]= -2045196100;
assign addr[52339]= -2067219829;
assign addr[52340]= -2086621133;
assign addr[52341]= -2103375398;
assign addr[52342]= -2117461370;
assign addr[52343]= -2128861181;
assign addr[52344]= -2137560369;
assign addr[52345]= -2143547897;
assign addr[52346]= -2146816171;
assign addr[52347]= -2147361045;
assign addr[52348]= -2145181827;
assign addr[52349]= -2140281282;
assign addr[52350]= -2132665626;
assign addr[52351]= -2122344521;
assign addr[52352]= -2109331059;
assign addr[52353]= -2093641749;
assign addr[52354]= -2075296495;
assign addr[52355]= -2054318569;
assign addr[52356]= -2030734582;
assign addr[52357]= -2004574453;
assign addr[52358]= -1975871368;
assign addr[52359]= -1944661739;
assign addr[52360]= -1910985158;
assign addr[52361]= -1874884346;
assign addr[52362]= -1836405100;
assign addr[52363]= -1795596234;
assign addr[52364]= -1752509516;
assign addr[52365]= -1707199606;
assign addr[52366]= -1659723983;
assign addr[52367]= -1610142873;
assign addr[52368]= -1558519173;
assign addr[52369]= -1504918373;
assign addr[52370]= -1449408469;
assign addr[52371]= -1392059879;
assign addr[52372]= -1332945355;
assign addr[52373]= -1272139887;
assign addr[52374]= -1209720613;
assign addr[52375]= -1145766716;
assign addr[52376]= -1080359326;
assign addr[52377]= -1013581418;
assign addr[52378]= -945517704;
assign addr[52379]= -876254528;
assign addr[52380]= -805879757;
assign addr[52381]= -734482665;
assign addr[52382]= -662153826;
assign addr[52383]= -588984994;
assign addr[52384]= -515068990;
assign addr[52385]= -440499581;
assign addr[52386]= -365371365;
assign addr[52387]= -289779648;
assign addr[52388]= -213820322;
assign addr[52389]= -137589750;
assign addr[52390]= -61184634;
assign addr[52391]= 15298099;
assign addr[52392]= 91761426;
assign addr[52393]= 168108346;
assign addr[52394]= 244242007;
assign addr[52395]= 320065829;
assign addr[52396]= 395483624;
assign addr[52397]= 470399716;
assign addr[52398]= 544719071;
assign addr[52399]= 618347408;
assign addr[52400]= 691191324;
assign addr[52401]= 763158411;
assign addr[52402]= 834157373;
assign addr[52403]= 904098143;
assign addr[52404]= 972891995;
assign addr[52405]= 1040451659;
assign addr[52406]= 1106691431;
assign addr[52407]= 1171527280;
assign addr[52408]= 1234876957;
assign addr[52409]= 1296660098;
assign addr[52410]= 1356798326;
assign addr[52411]= 1415215352;
assign addr[52412]= 1471837070;
assign addr[52413]= 1526591649;
assign addr[52414]= 1579409630;
assign addr[52415]= 1630224009;
assign addr[52416]= 1678970324;
assign addr[52417]= 1725586737;
assign addr[52418]= 1770014111;
assign addr[52419]= 1812196087;
assign addr[52420]= 1852079154;
assign addr[52421]= 1889612716;
assign addr[52422]= 1924749160;
assign addr[52423]= 1957443913;
assign addr[52424]= 1987655498;
assign addr[52425]= 2015345591;
assign addr[52426]= 2040479063;
assign addr[52427]= 2063024031;
assign addr[52428]= 2082951896;
assign addr[52429]= 2100237377;
assign addr[52430]= 2114858546;
assign addr[52431]= 2126796855;
assign addr[52432]= 2136037160;
assign addr[52433]= 2142567738;
assign addr[52434]= 2146380306;
assign addr[52435]= 2147470025;
assign addr[52436]= 2145835515;
assign addr[52437]= 2141478848;
assign addr[52438]= 2134405552;
assign addr[52439]= 2124624598;
assign addr[52440]= 2112148396;
assign addr[52441]= 2096992772;
assign addr[52442]= 2079176953;
assign addr[52443]= 2058723538;
assign addr[52444]= 2035658475;
assign addr[52445]= 2010011024;
assign addr[52446]= 1981813720;
assign addr[52447]= 1951102334;
assign addr[52448]= 1917915825;
assign addr[52449]= 1882296293;
assign addr[52450]= 1844288924;
assign addr[52451]= 1803941934;
assign addr[52452]= 1761306505;
assign addr[52453]= 1716436725;
assign addr[52454]= 1669389513;
assign addr[52455]= 1620224553;
assign addr[52456]= 1569004214;
assign addr[52457]= 1515793473;
assign addr[52458]= 1460659832;
assign addr[52459]= 1403673233;
assign addr[52460]= 1344905966;
assign addr[52461]= 1284432584;
assign addr[52462]= 1222329801;
assign addr[52463]= 1158676398;
assign addr[52464]= 1093553126;
assign addr[52465]= 1027042599;
assign addr[52466]= 959229189;
assign addr[52467]= 890198924;
assign addr[52468]= 820039373;
assign addr[52469]= 748839539;
assign addr[52470]= 676689746;
assign addr[52471]= 603681519;
assign addr[52472]= 529907477;
assign addr[52473]= 455461206;
assign addr[52474]= 380437148;
assign addr[52475]= 304930476;
assign addr[52476]= 229036977;
assign addr[52477]= 152852926;
assign addr[52478]= 76474970;
assign addr[52479]= 0;
assign addr[52480]= -76474970;
assign addr[52481]= -152852926;
assign addr[52482]= -229036977;
assign addr[52483]= -304930476;
assign addr[52484]= -380437148;
assign addr[52485]= -455461206;
assign addr[52486]= -529907477;
assign addr[52487]= -603681519;
assign addr[52488]= -676689746;
assign addr[52489]= -748839539;
assign addr[52490]= -820039373;
assign addr[52491]= -890198924;
assign addr[52492]= -959229189;
assign addr[52493]= -1027042599;
assign addr[52494]= -1093553126;
assign addr[52495]= -1158676398;
assign addr[52496]= -1222329801;
assign addr[52497]= -1284432584;
assign addr[52498]= -1344905966;
assign addr[52499]= -1403673233;
assign addr[52500]= -1460659832;
assign addr[52501]= -1515793473;
assign addr[52502]= -1569004214;
assign addr[52503]= -1620224553;
assign addr[52504]= -1669389513;
assign addr[52505]= -1716436725;
assign addr[52506]= -1761306505;
assign addr[52507]= -1803941934;
assign addr[52508]= -1844288924;
assign addr[52509]= -1882296293;
assign addr[52510]= -1917915825;
assign addr[52511]= -1951102334;
assign addr[52512]= -1981813720;
assign addr[52513]= -2010011024;
assign addr[52514]= -2035658475;
assign addr[52515]= -2058723538;
assign addr[52516]= -2079176953;
assign addr[52517]= -2096992772;
assign addr[52518]= -2112148396;
assign addr[52519]= -2124624598;
assign addr[52520]= -2134405552;
assign addr[52521]= -2141478848;
assign addr[52522]= -2145835515;
assign addr[52523]= -2147470025;
assign addr[52524]= -2146380306;
assign addr[52525]= -2142567738;
assign addr[52526]= -2136037160;
assign addr[52527]= -2126796855;
assign addr[52528]= -2114858546;
assign addr[52529]= -2100237377;
assign addr[52530]= -2082951896;
assign addr[52531]= -2063024031;
assign addr[52532]= -2040479063;
assign addr[52533]= -2015345591;
assign addr[52534]= -1987655498;
assign addr[52535]= -1957443913;
assign addr[52536]= -1924749160;
assign addr[52537]= -1889612716;
assign addr[52538]= -1852079154;
assign addr[52539]= -1812196087;
assign addr[52540]= -1770014111;
assign addr[52541]= -1725586737;
assign addr[52542]= -1678970324;
assign addr[52543]= -1630224009;
assign addr[52544]= -1579409630;
assign addr[52545]= -1526591649;
assign addr[52546]= -1471837070;
assign addr[52547]= -1415215352;
assign addr[52548]= -1356798326;
assign addr[52549]= -1296660098;
assign addr[52550]= -1234876957;
assign addr[52551]= -1171527280;
assign addr[52552]= -1106691431;
assign addr[52553]= -1040451659;
assign addr[52554]= -972891995;
assign addr[52555]= -904098143;
assign addr[52556]= -834157373;
assign addr[52557]= -763158411;
assign addr[52558]= -691191324;
assign addr[52559]= -618347408;
assign addr[52560]= -544719071;
assign addr[52561]= -470399716;
assign addr[52562]= -395483624;
assign addr[52563]= -320065829;
assign addr[52564]= -244242007;
assign addr[52565]= -168108346;
assign addr[52566]= -91761426;
assign addr[52567]= -15298099;
assign addr[52568]= 61184634;
assign addr[52569]= 137589750;
assign addr[52570]= 213820322;
assign addr[52571]= 289779648;
assign addr[52572]= 365371365;
assign addr[52573]= 440499581;
assign addr[52574]= 515068990;
assign addr[52575]= 588984994;
assign addr[52576]= 662153826;
assign addr[52577]= 734482665;
assign addr[52578]= 805879757;
assign addr[52579]= 876254528;
assign addr[52580]= 945517704;
assign addr[52581]= 1013581418;
assign addr[52582]= 1080359326;
assign addr[52583]= 1145766716;
assign addr[52584]= 1209720613;
assign addr[52585]= 1272139887;
assign addr[52586]= 1332945355;
assign addr[52587]= 1392059879;
assign addr[52588]= 1449408469;
assign addr[52589]= 1504918373;
assign addr[52590]= 1558519173;
assign addr[52591]= 1610142873;
assign addr[52592]= 1659723983;
assign addr[52593]= 1707199606;
assign addr[52594]= 1752509516;
assign addr[52595]= 1795596234;
assign addr[52596]= 1836405100;
assign addr[52597]= 1874884346;
assign addr[52598]= 1910985158;
assign addr[52599]= 1944661739;
assign addr[52600]= 1975871368;
assign addr[52601]= 2004574453;
assign addr[52602]= 2030734582;
assign addr[52603]= 2054318569;
assign addr[52604]= 2075296495;
assign addr[52605]= 2093641749;
assign addr[52606]= 2109331059;
assign addr[52607]= 2122344521;
assign addr[52608]= 2132665626;
assign addr[52609]= 2140281282;
assign addr[52610]= 2145181827;
assign addr[52611]= 2147361045;
assign addr[52612]= 2146816171;
assign addr[52613]= 2143547897;
assign addr[52614]= 2137560369;
assign addr[52615]= 2128861181;
assign addr[52616]= 2117461370;
assign addr[52617]= 2103375398;
assign addr[52618]= 2086621133;
assign addr[52619]= 2067219829;
assign addr[52620]= 2045196100;
assign addr[52621]= 2020577882;
assign addr[52622]= 1993396407;
assign addr[52623]= 1963686155;
assign addr[52624]= 1931484818;
assign addr[52625]= 1896833245;
assign addr[52626]= 1859775393;
assign addr[52627]= 1820358275;
assign addr[52628]= 1778631892;
assign addr[52629]= 1734649179;
assign addr[52630]= 1688465931;
assign addr[52631]= 1640140734;
assign addr[52632]= 1589734894;
assign addr[52633]= 1537312353;
assign addr[52634]= 1482939614;
assign addr[52635]= 1426685652;
assign addr[52636]= 1368621831;
assign addr[52637]= 1308821808;
assign addr[52638]= 1247361445;
assign addr[52639]= 1184318708;
assign addr[52640]= 1119773573;
assign addr[52641]= 1053807919;
assign addr[52642]= 986505429;
assign addr[52643]= 917951481;
assign addr[52644]= 848233042;
assign addr[52645]= 777438554;
assign addr[52646]= 705657826;
assign addr[52647]= 632981917;
assign addr[52648]= 559503022;
assign addr[52649]= 485314355;
assign addr[52650]= 410510029;
assign addr[52651]= 335184940;
assign addr[52652]= 259434643;
assign addr[52653]= 183355234;
assign addr[52654]= 107043224;
assign addr[52655]= 30595422;
assign addr[52656]= -45891193;
assign addr[52657]= -122319591;
assign addr[52658]= -198592817;
assign addr[52659]= -274614114;
assign addr[52660]= -350287041;
assign addr[52661]= -425515602;
assign addr[52662]= -500204365;
assign addr[52663]= -574258580;
assign addr[52664]= -647584304;
assign addr[52665]= -720088517;
assign addr[52666]= -791679244;
assign addr[52667]= -862265664;
assign addr[52668]= -931758235;
assign addr[52669]= -1000068799;
assign addr[52670]= -1067110699;
assign addr[52671]= -1132798888;
assign addr[52672]= -1197050035;
assign addr[52673]= -1259782632;
assign addr[52674]= -1320917099;
assign addr[52675]= -1380375881;
assign addr[52676]= -1438083551;
assign addr[52677]= -1493966902;
assign addr[52678]= -1547955041;
assign addr[52679]= -1599979481;
assign addr[52680]= -1649974225;
assign addr[52681]= -1697875851;
assign addr[52682]= -1743623590;
assign addr[52683]= -1787159411;
assign addr[52684]= -1828428082;
assign addr[52685]= -1867377253;
assign addr[52686]= -1903957513;
assign addr[52687]= -1938122457;
assign addr[52688]= -1969828744;
assign addr[52689]= -1999036154;
assign addr[52690]= -2025707632;
assign addr[52691]= -2049809346;
assign addr[52692]= -2071310720;
assign addr[52693]= -2090184478;
assign addr[52694]= -2106406677;
assign addr[52695]= -2119956737;
assign addr[52696]= -2130817471;
assign addr[52697]= -2138975100;
assign addr[52698]= -2144419275;
assign addr[52699]= -2147143090;
assign addr[52700]= -2147143090;
assign addr[52701]= -2144419275;
assign addr[52702]= -2138975100;
assign addr[52703]= -2130817471;
assign addr[52704]= -2119956737;
assign addr[52705]= -2106406677;
assign addr[52706]= -2090184478;
assign addr[52707]= -2071310720;
assign addr[52708]= -2049809346;
assign addr[52709]= -2025707632;
assign addr[52710]= -1999036154;
assign addr[52711]= -1969828744;
assign addr[52712]= -1938122457;
assign addr[52713]= -1903957513;
assign addr[52714]= -1867377253;
assign addr[52715]= -1828428082;
assign addr[52716]= -1787159411;
assign addr[52717]= -1743623590;
assign addr[52718]= -1697875851;
assign addr[52719]= -1649974225;
assign addr[52720]= -1599979481;
assign addr[52721]= -1547955041;
assign addr[52722]= -1493966902;
assign addr[52723]= -1438083551;
assign addr[52724]= -1380375881;
assign addr[52725]= -1320917099;
assign addr[52726]= -1259782632;
assign addr[52727]= -1197050035;
assign addr[52728]= -1132798888;
assign addr[52729]= -1067110699;
assign addr[52730]= -1000068799;
assign addr[52731]= -931758235;
assign addr[52732]= -862265664;
assign addr[52733]= -791679244;
assign addr[52734]= -720088517;
assign addr[52735]= -647584304;
assign addr[52736]= -574258580;
assign addr[52737]= -500204365;
assign addr[52738]= -425515602;
assign addr[52739]= -350287041;
assign addr[52740]= -274614114;
assign addr[52741]= -198592817;
assign addr[52742]= -122319591;
assign addr[52743]= -45891193;
assign addr[52744]= 30595422;
assign addr[52745]= 107043224;
assign addr[52746]= 183355234;
assign addr[52747]= 259434643;
assign addr[52748]= 335184940;
assign addr[52749]= 410510029;
assign addr[52750]= 485314355;
assign addr[52751]= 559503022;
assign addr[52752]= 632981917;
assign addr[52753]= 705657826;
assign addr[52754]= 777438554;
assign addr[52755]= 848233042;
assign addr[52756]= 917951481;
assign addr[52757]= 986505429;
assign addr[52758]= 1053807919;
assign addr[52759]= 1119773573;
assign addr[52760]= 1184318708;
assign addr[52761]= 1247361445;
assign addr[52762]= 1308821808;
assign addr[52763]= 1368621831;
assign addr[52764]= 1426685652;
assign addr[52765]= 1482939614;
assign addr[52766]= 1537312353;
assign addr[52767]= 1589734894;
assign addr[52768]= 1640140734;
assign addr[52769]= 1688465931;
assign addr[52770]= 1734649179;
assign addr[52771]= 1778631892;
assign addr[52772]= 1820358275;
assign addr[52773]= 1859775393;
assign addr[52774]= 1896833245;
assign addr[52775]= 1931484818;
assign addr[52776]= 1963686155;
assign addr[52777]= 1993396407;
assign addr[52778]= 2020577882;
assign addr[52779]= 2045196100;
assign addr[52780]= 2067219829;
assign addr[52781]= 2086621133;
assign addr[52782]= 2103375398;
assign addr[52783]= 2117461370;
assign addr[52784]= 2128861181;
assign addr[52785]= 2137560369;
assign addr[52786]= 2143547897;
assign addr[52787]= 2146816171;
assign addr[52788]= 2147361045;
assign addr[52789]= 2145181827;
assign addr[52790]= 2140281282;
assign addr[52791]= 2132665626;
assign addr[52792]= 2122344521;
assign addr[52793]= 2109331059;
assign addr[52794]= 2093641749;
assign addr[52795]= 2075296495;
assign addr[52796]= 2054318569;
assign addr[52797]= 2030734582;
assign addr[52798]= 2004574453;
assign addr[52799]= 1975871368;
assign addr[52800]= 1944661739;
assign addr[52801]= 1910985158;
assign addr[52802]= 1874884346;
assign addr[52803]= 1836405100;
assign addr[52804]= 1795596234;
assign addr[52805]= 1752509516;
assign addr[52806]= 1707199606;
assign addr[52807]= 1659723983;
assign addr[52808]= 1610142873;
assign addr[52809]= 1558519173;
assign addr[52810]= 1504918373;
assign addr[52811]= 1449408469;
assign addr[52812]= 1392059879;
assign addr[52813]= 1332945355;
assign addr[52814]= 1272139887;
assign addr[52815]= 1209720613;
assign addr[52816]= 1145766716;
assign addr[52817]= 1080359326;
assign addr[52818]= 1013581418;
assign addr[52819]= 945517704;
assign addr[52820]= 876254528;
assign addr[52821]= 805879757;
assign addr[52822]= 734482665;
assign addr[52823]= 662153826;
assign addr[52824]= 588984994;
assign addr[52825]= 515068990;
assign addr[52826]= 440499581;
assign addr[52827]= 365371365;
assign addr[52828]= 289779648;
assign addr[52829]= 213820322;
assign addr[52830]= 137589750;
assign addr[52831]= 61184634;
assign addr[52832]= -15298099;
assign addr[52833]= -91761426;
assign addr[52834]= -168108346;
assign addr[52835]= -244242007;
assign addr[52836]= -320065829;
assign addr[52837]= -395483624;
assign addr[52838]= -470399716;
assign addr[52839]= -544719071;
assign addr[52840]= -618347408;
assign addr[52841]= -691191324;
assign addr[52842]= -763158411;
assign addr[52843]= -834157373;
assign addr[52844]= -904098143;
assign addr[52845]= -972891995;
assign addr[52846]= -1040451659;
assign addr[52847]= -1106691431;
assign addr[52848]= -1171527280;
assign addr[52849]= -1234876957;
assign addr[52850]= -1296660098;
assign addr[52851]= -1356798326;
assign addr[52852]= -1415215352;
assign addr[52853]= -1471837070;
assign addr[52854]= -1526591649;
assign addr[52855]= -1579409630;
assign addr[52856]= -1630224009;
assign addr[52857]= -1678970324;
assign addr[52858]= -1725586737;
assign addr[52859]= -1770014111;
assign addr[52860]= -1812196087;
assign addr[52861]= -1852079154;
assign addr[52862]= -1889612716;
assign addr[52863]= -1924749160;
assign addr[52864]= -1957443913;
assign addr[52865]= -1987655498;
assign addr[52866]= -2015345591;
assign addr[52867]= -2040479063;
assign addr[52868]= -2063024031;
assign addr[52869]= -2082951896;
assign addr[52870]= -2100237377;
assign addr[52871]= -2114858546;
assign addr[52872]= -2126796855;
assign addr[52873]= -2136037160;
assign addr[52874]= -2142567738;
assign addr[52875]= -2146380306;
assign addr[52876]= -2147470025;
assign addr[52877]= -2145835515;
assign addr[52878]= -2141478848;
assign addr[52879]= -2134405552;
assign addr[52880]= -2124624598;
assign addr[52881]= -2112148396;
assign addr[52882]= -2096992772;
assign addr[52883]= -2079176953;
assign addr[52884]= -2058723538;
assign addr[52885]= -2035658475;
assign addr[52886]= -2010011024;
assign addr[52887]= -1981813720;
assign addr[52888]= -1951102334;
assign addr[52889]= -1917915825;
assign addr[52890]= -1882296293;
assign addr[52891]= -1844288924;
assign addr[52892]= -1803941934;
assign addr[52893]= -1761306505;
assign addr[52894]= -1716436725;
assign addr[52895]= -1669389513;
assign addr[52896]= -1620224553;
assign addr[52897]= -1569004214;
assign addr[52898]= -1515793473;
assign addr[52899]= -1460659832;
assign addr[52900]= -1403673233;
assign addr[52901]= -1344905966;
assign addr[52902]= -1284432584;
assign addr[52903]= -1222329801;
assign addr[52904]= -1158676398;
assign addr[52905]= -1093553126;
assign addr[52906]= -1027042599;
assign addr[52907]= -959229189;
assign addr[52908]= -890198924;
assign addr[52909]= -820039373;
assign addr[52910]= -748839539;
assign addr[52911]= -676689746;
assign addr[52912]= -603681519;
assign addr[52913]= -529907477;
assign addr[52914]= -455461206;
assign addr[52915]= -380437148;
assign addr[52916]= -304930476;
assign addr[52917]= -229036977;
assign addr[52918]= -152852926;
assign addr[52919]= -76474970;
assign addr[52920]= 0;
assign addr[52921]= 76474970;
assign addr[52922]= 152852926;
assign addr[52923]= 229036977;
assign addr[52924]= 304930476;
assign addr[52925]= 380437148;
assign addr[52926]= 455461206;
assign addr[52927]= 529907477;
assign addr[52928]= 603681519;
assign addr[52929]= 676689746;
assign addr[52930]= 748839539;
assign addr[52931]= 820039373;
assign addr[52932]= 890198924;
assign addr[52933]= 959229189;
assign addr[52934]= 1027042599;
assign addr[52935]= 1093553126;
assign addr[52936]= 1158676398;
assign addr[52937]= 1222329801;
assign addr[52938]= 1284432584;
assign addr[52939]= 1344905966;
assign addr[52940]= 1403673233;
assign addr[52941]= 1460659832;
assign addr[52942]= 1515793473;
assign addr[52943]= 1569004214;
assign addr[52944]= 1620224553;
assign addr[52945]= 1669389513;
assign addr[52946]= 1716436725;
assign addr[52947]= 1761306505;
assign addr[52948]= 1803941934;
assign addr[52949]= 1844288924;
assign addr[52950]= 1882296293;
assign addr[52951]= 1917915825;
assign addr[52952]= 1951102334;
assign addr[52953]= 1981813720;
assign addr[52954]= 2010011024;
assign addr[52955]= 2035658475;
assign addr[52956]= 2058723538;
assign addr[52957]= 2079176953;
assign addr[52958]= 2096992772;
assign addr[52959]= 2112148396;
assign addr[52960]= 2124624598;
assign addr[52961]= 2134405552;
assign addr[52962]= 2141478848;
assign addr[52963]= 2145835515;
assign addr[52964]= 2147470025;
assign addr[52965]= 2146380306;
assign addr[52966]= 2142567738;
assign addr[52967]= 2136037160;
assign addr[52968]= 2126796855;
assign addr[52969]= 2114858546;
assign addr[52970]= 2100237377;
assign addr[52971]= 2082951896;
assign addr[52972]= 2063024031;
assign addr[52973]= 2040479063;
assign addr[52974]= 2015345591;
assign addr[52975]= 1987655498;
assign addr[52976]= 1957443913;
assign addr[52977]= 1924749160;
assign addr[52978]= 1889612716;
assign addr[52979]= 1852079154;
assign addr[52980]= 1812196087;
assign addr[52981]= 1770014111;
assign addr[52982]= 1725586737;
assign addr[52983]= 1678970324;
assign addr[52984]= 1630224009;
assign addr[52985]= 1579409630;
assign addr[52986]= 1526591649;
assign addr[52987]= 1471837070;
assign addr[52988]= 1415215352;
assign addr[52989]= 1356798326;
assign addr[52990]= 1296660098;
assign addr[52991]= 1234876957;
assign addr[52992]= 1171527280;
assign addr[52993]= 1106691431;
assign addr[52994]= 1040451659;
assign addr[52995]= 972891995;
assign addr[52996]= 904098143;
assign addr[52997]= 834157373;
assign addr[52998]= 763158411;
assign addr[52999]= 691191324;
assign addr[53000]= 618347408;
assign addr[53001]= 544719071;
assign addr[53002]= 470399716;
assign addr[53003]= 395483624;
assign addr[53004]= 320065829;
assign addr[53005]= 244242007;
assign addr[53006]= 168108346;
assign addr[53007]= 91761426;
assign addr[53008]= 15298099;
assign addr[53009]= -61184634;
assign addr[53010]= -137589750;
assign addr[53011]= -213820322;
assign addr[53012]= -289779648;
assign addr[53013]= -365371365;
assign addr[53014]= -440499581;
assign addr[53015]= -515068990;
assign addr[53016]= -588984994;
assign addr[53017]= -662153826;
assign addr[53018]= -734482665;
assign addr[53019]= -805879757;
assign addr[53020]= -876254528;
assign addr[53021]= -945517704;
assign addr[53022]= -1013581418;
assign addr[53023]= -1080359326;
assign addr[53024]= -1145766716;
assign addr[53025]= -1209720613;
assign addr[53026]= -1272139887;
assign addr[53027]= -1332945355;
assign addr[53028]= -1392059879;
assign addr[53029]= -1449408469;
assign addr[53030]= -1504918373;
assign addr[53031]= -1558519173;
assign addr[53032]= -1610142873;
assign addr[53033]= -1659723983;
assign addr[53034]= -1707199606;
assign addr[53035]= -1752509516;
assign addr[53036]= -1795596234;
assign addr[53037]= -1836405100;
assign addr[53038]= -1874884346;
assign addr[53039]= -1910985158;
assign addr[53040]= -1944661739;
assign addr[53041]= -1975871368;
assign addr[53042]= -2004574453;
assign addr[53043]= -2030734582;
assign addr[53044]= -2054318569;
assign addr[53045]= -2075296495;
assign addr[53046]= -2093641749;
assign addr[53047]= -2109331059;
assign addr[53048]= -2122344521;
assign addr[53049]= -2132665626;
assign addr[53050]= -2140281282;
assign addr[53051]= -2145181827;
assign addr[53052]= -2147361045;
assign addr[53053]= -2146816171;
assign addr[53054]= -2143547897;
assign addr[53055]= -2137560369;
assign addr[53056]= -2128861181;
assign addr[53057]= -2117461370;
assign addr[53058]= -2103375398;
assign addr[53059]= -2086621133;
assign addr[53060]= -2067219829;
assign addr[53061]= -2045196100;
assign addr[53062]= -2020577882;
assign addr[53063]= -1993396407;
assign addr[53064]= -1963686155;
assign addr[53065]= -1931484818;
assign addr[53066]= -1896833245;
assign addr[53067]= -1859775393;
assign addr[53068]= -1820358275;
assign addr[53069]= -1778631892;
assign addr[53070]= -1734649179;
assign addr[53071]= -1688465931;
assign addr[53072]= -1640140734;
assign addr[53073]= -1589734894;
assign addr[53074]= -1537312353;
assign addr[53075]= -1482939614;
assign addr[53076]= -1426685652;
assign addr[53077]= -1368621831;
assign addr[53078]= -1308821808;
assign addr[53079]= -1247361445;
assign addr[53080]= -1184318708;
assign addr[53081]= -1119773573;
assign addr[53082]= -1053807919;
assign addr[53083]= -986505429;
assign addr[53084]= -917951481;
assign addr[53085]= -848233042;
assign addr[53086]= -777438554;
assign addr[53087]= -705657826;
assign addr[53088]= -632981917;
assign addr[53089]= -559503022;
assign addr[53090]= -485314355;
assign addr[53091]= -410510029;
assign addr[53092]= -335184940;
assign addr[53093]= -259434643;
assign addr[53094]= -183355234;
assign addr[53095]= -107043224;
assign addr[53096]= -30595422;
assign addr[53097]= 45891193;
assign addr[53098]= 122319591;
assign addr[53099]= 198592817;
assign addr[53100]= 274614114;
assign addr[53101]= 350287041;
assign addr[53102]= 425515602;
assign addr[53103]= 500204365;
assign addr[53104]= 574258580;
assign addr[53105]= 647584304;
assign addr[53106]= 720088517;
assign addr[53107]= 791679244;
assign addr[53108]= 862265664;
assign addr[53109]= 931758235;
assign addr[53110]= 1000068799;
assign addr[53111]= 1067110699;
assign addr[53112]= 1132798888;
assign addr[53113]= 1197050035;
assign addr[53114]= 1259782632;
assign addr[53115]= 1320917099;
assign addr[53116]= 1380375881;
assign addr[53117]= 1438083551;
assign addr[53118]= 1493966902;
assign addr[53119]= 1547955041;
assign addr[53120]= 1599979481;
assign addr[53121]= 1649974225;
assign addr[53122]= 1697875851;
assign addr[53123]= 1743623590;
assign addr[53124]= 1787159411;
assign addr[53125]= 1828428082;
assign addr[53126]= 1867377253;
assign addr[53127]= 1903957513;
assign addr[53128]= 1938122457;
assign addr[53129]= 1969828744;
assign addr[53130]= 1999036154;
assign addr[53131]= 2025707632;
assign addr[53132]= 2049809346;
assign addr[53133]= 2071310720;
assign addr[53134]= 2090184478;
assign addr[53135]= 2106406677;
assign addr[53136]= 2119956737;
assign addr[53137]= 2130817471;
assign addr[53138]= 2138975100;
assign addr[53139]= 2144419275;
assign addr[53140]= 2147143090;
assign addr[53141]= 2147143090;
assign addr[53142]= 2144419275;
assign addr[53143]= 2138975100;
assign addr[53144]= 2130817471;
assign addr[53145]= 2119956737;
assign addr[53146]= 2106406677;
assign addr[53147]= 2090184478;
assign addr[53148]= 2071310720;
assign addr[53149]= 2049809346;
assign addr[53150]= 2025707632;
assign addr[53151]= 1999036154;
assign addr[53152]= 1969828744;
assign addr[53153]= 1938122457;
assign addr[53154]= 1903957513;
assign addr[53155]= 1867377253;
assign addr[53156]= 1828428082;
assign addr[53157]= 1787159411;
assign addr[53158]= 1743623590;
assign addr[53159]= 1697875851;
assign addr[53160]= 1649974225;
assign addr[53161]= 1599979481;
assign addr[53162]= 1547955041;
assign addr[53163]= 1493966902;
assign addr[53164]= 1438083551;
assign addr[53165]= 1380375881;
assign addr[53166]= 1320917099;
assign addr[53167]= 1259782632;
assign addr[53168]= 1197050035;
assign addr[53169]= 1132798888;
assign addr[53170]= 1067110699;
assign addr[53171]= 1000068799;
assign addr[53172]= 931758235;
assign addr[53173]= 862265664;
assign addr[53174]= 791679244;
assign addr[53175]= 720088517;
assign addr[53176]= 647584304;
assign addr[53177]= 574258580;
assign addr[53178]= 500204365;
assign addr[53179]= 425515602;
assign addr[53180]= 350287041;
assign addr[53181]= 274614114;
assign addr[53182]= 198592817;
assign addr[53183]= 122319591;
assign addr[53184]= 45891193;
assign addr[53185]= -30595422;
assign addr[53186]= -107043224;
assign addr[53187]= -183355234;
assign addr[53188]= -259434643;
assign addr[53189]= -335184940;
assign addr[53190]= -410510029;
assign addr[53191]= -485314355;
assign addr[53192]= -559503022;
assign addr[53193]= -632981917;
assign addr[53194]= -705657826;
assign addr[53195]= -777438554;
assign addr[53196]= -848233042;
assign addr[53197]= -917951481;
assign addr[53198]= -986505429;
assign addr[53199]= -1053807919;
assign addr[53200]= -1119773573;
assign addr[53201]= -1184318708;
assign addr[53202]= -1247361445;
assign addr[53203]= -1308821808;
assign addr[53204]= -1368621831;
assign addr[53205]= -1426685652;
assign addr[53206]= -1482939614;
assign addr[53207]= -1537312353;
assign addr[53208]= -1589734894;
assign addr[53209]= -1640140734;
assign addr[53210]= -1688465931;
assign addr[53211]= -1734649179;
assign addr[53212]= -1778631892;
assign addr[53213]= -1820358275;
assign addr[53214]= -1859775393;
assign addr[53215]= -1896833245;
assign addr[53216]= -1931484818;
assign addr[53217]= -1963686155;
assign addr[53218]= -1993396407;
assign addr[53219]= -2020577882;
assign addr[53220]= -2045196100;
assign addr[53221]= -2067219829;
assign addr[53222]= -2086621133;
assign addr[53223]= -2103375398;
assign addr[53224]= -2117461370;
assign addr[53225]= -2128861181;
assign addr[53226]= -2137560369;
assign addr[53227]= -2143547897;
assign addr[53228]= -2146816171;
assign addr[53229]= -2147361045;
assign addr[53230]= -2145181827;
assign addr[53231]= -2140281282;
assign addr[53232]= -2132665626;
assign addr[53233]= -2122344521;
assign addr[53234]= -2109331059;
assign addr[53235]= -2093641749;
assign addr[53236]= -2075296495;
assign addr[53237]= -2054318569;
assign addr[53238]= -2030734582;
assign addr[53239]= -2004574453;
assign addr[53240]= -1975871368;
assign addr[53241]= -1944661739;
assign addr[53242]= -1910985158;
assign addr[53243]= -1874884346;
assign addr[53244]= -1836405100;
assign addr[53245]= -1795596234;
assign addr[53246]= -1752509516;
assign addr[53247]= -1707199606;
assign addr[53248]= -1659723983;
assign addr[53249]= -1610142873;
assign addr[53250]= -1558519173;
assign addr[53251]= -1504918373;
assign addr[53252]= -1449408469;
assign addr[53253]= -1392059879;
assign addr[53254]= -1332945355;
assign addr[53255]= -1272139887;
assign addr[53256]= -1209720613;
assign addr[53257]= -1145766716;
assign addr[53258]= -1080359326;
assign addr[53259]= -1013581418;
assign addr[53260]= -945517704;
assign addr[53261]= -876254528;
assign addr[53262]= -805879757;
assign addr[53263]= -734482665;
assign addr[53264]= -662153826;
assign addr[53265]= -588984994;
assign addr[53266]= -515068990;
assign addr[53267]= -440499581;
assign addr[53268]= -365371365;
assign addr[53269]= -289779648;
assign addr[53270]= -213820322;
assign addr[53271]= -137589750;
assign addr[53272]= -61184634;
assign addr[53273]= 15298099;
assign addr[53274]= 91761426;
assign addr[53275]= 168108346;
assign addr[53276]= 244242007;
assign addr[53277]= 320065829;
assign addr[53278]= 395483624;
assign addr[53279]= 470399716;
assign addr[53280]= 544719071;
assign addr[53281]= 618347408;
assign addr[53282]= 691191324;
assign addr[53283]= 763158411;
assign addr[53284]= 834157373;
assign addr[53285]= 904098143;
assign addr[53286]= 972891995;
assign addr[53287]= 1040451659;
assign addr[53288]= 1106691431;
assign addr[53289]= 1171527280;
assign addr[53290]= 1234876957;
assign addr[53291]= 1296660098;
assign addr[53292]= 1356798326;
assign addr[53293]= 1415215352;
assign addr[53294]= 1471837070;
assign addr[53295]= 1526591649;
assign addr[53296]= 1579409630;
assign addr[53297]= 1630224009;
assign addr[53298]= 1678970324;
assign addr[53299]= 1725586737;
assign addr[53300]= 1770014111;
assign addr[53301]= 1812196087;
assign addr[53302]= 1852079154;
assign addr[53303]= 1889612716;
assign addr[53304]= 1924749160;
assign addr[53305]= 1957443913;
assign addr[53306]= 1987655498;
assign addr[53307]= 2015345591;
assign addr[53308]= 2040479063;
assign addr[53309]= 2063024031;
assign addr[53310]= 2082951896;
assign addr[53311]= 2100237377;
assign addr[53312]= 2114858546;
assign addr[53313]= 2126796855;
assign addr[53314]= 2136037160;
assign addr[53315]= 2142567738;
assign addr[53316]= 2146380306;
assign addr[53317]= 2147470025;
assign addr[53318]= 2145835515;
assign addr[53319]= 2141478848;
assign addr[53320]= 2134405552;
assign addr[53321]= 2124624598;
assign addr[53322]= 2112148396;
assign addr[53323]= 2096992772;
assign addr[53324]= 2079176953;
assign addr[53325]= 2058723538;
assign addr[53326]= 2035658475;
assign addr[53327]= 2010011024;
assign addr[53328]= 1981813720;
assign addr[53329]= 1951102334;
assign addr[53330]= 1917915825;
assign addr[53331]= 1882296293;
assign addr[53332]= 1844288924;
assign addr[53333]= 1803941934;
assign addr[53334]= 1761306505;
assign addr[53335]= 1716436725;
assign addr[53336]= 1669389513;
assign addr[53337]= 1620224553;
assign addr[53338]= 1569004214;
assign addr[53339]= 1515793473;
assign addr[53340]= 1460659832;
assign addr[53341]= 1403673233;
assign addr[53342]= 1344905966;
assign addr[53343]= 1284432584;
assign addr[53344]= 1222329801;
assign addr[53345]= 1158676398;
assign addr[53346]= 1093553126;
assign addr[53347]= 1027042599;
assign addr[53348]= 959229189;
assign addr[53349]= 890198924;
assign addr[53350]= 820039373;
assign addr[53351]= 748839539;
assign addr[53352]= 676689746;
assign addr[53353]= 603681519;
assign addr[53354]= 529907477;
assign addr[53355]= 455461206;
assign addr[53356]= 380437148;
assign addr[53357]= 304930476;
assign addr[53358]= 229036977;
assign addr[53359]= 152852926;
assign addr[53360]= 76474970;
assign addr[53361]= 0;
assign addr[53362]= -76474970;
assign addr[53363]= -152852926;
assign addr[53364]= -229036977;
assign addr[53365]= -304930476;
assign addr[53366]= -380437148;
assign addr[53367]= -455461206;
assign addr[53368]= -529907477;
assign addr[53369]= -603681519;
assign addr[53370]= -676689746;
assign addr[53371]= -748839539;
assign addr[53372]= -820039373;
assign addr[53373]= -890198924;
assign addr[53374]= -959229189;
assign addr[53375]= -1027042599;
assign addr[53376]= -1093553126;
assign addr[53377]= -1158676398;
assign addr[53378]= -1222329801;
assign addr[53379]= -1284432584;
assign addr[53380]= -1344905966;
assign addr[53381]= -1403673233;
assign addr[53382]= -1460659832;
assign addr[53383]= -1515793473;
assign addr[53384]= -1569004214;
assign addr[53385]= -1620224553;
assign addr[53386]= -1669389513;
assign addr[53387]= -1716436725;
assign addr[53388]= -1761306505;
assign addr[53389]= -1803941934;
assign addr[53390]= -1844288924;
assign addr[53391]= -1882296293;
assign addr[53392]= -1917915825;
assign addr[53393]= -1951102334;
assign addr[53394]= -1981813720;
assign addr[53395]= -2010011024;
assign addr[53396]= -2035658475;
assign addr[53397]= -2058723538;
assign addr[53398]= -2079176953;
assign addr[53399]= -2096992772;
assign addr[53400]= -2112148396;
assign addr[53401]= -2124624598;
assign addr[53402]= -2134405552;
assign addr[53403]= -2141478848;
assign addr[53404]= -2145835515;
assign addr[53405]= -2147470025;
assign addr[53406]= -2146380306;
assign addr[53407]= -2142567738;
assign addr[53408]= -2136037160;
assign addr[53409]= -2126796855;
assign addr[53410]= -2114858546;
assign addr[53411]= -2100237377;
assign addr[53412]= -2082951896;
assign addr[53413]= -2063024031;
assign addr[53414]= -2040479063;
assign addr[53415]= -2015345591;
assign addr[53416]= -1987655498;
assign addr[53417]= -1957443913;
assign addr[53418]= -1924749160;
assign addr[53419]= -1889612716;
assign addr[53420]= -1852079154;
assign addr[53421]= -1812196087;
assign addr[53422]= -1770014111;
assign addr[53423]= -1725586737;
assign addr[53424]= -1678970324;
assign addr[53425]= -1630224009;
assign addr[53426]= -1579409630;
assign addr[53427]= -1526591649;
assign addr[53428]= -1471837070;
assign addr[53429]= -1415215352;
assign addr[53430]= -1356798326;
assign addr[53431]= -1296660098;
assign addr[53432]= -1234876957;
assign addr[53433]= -1171527280;
assign addr[53434]= -1106691431;
assign addr[53435]= -1040451659;
assign addr[53436]= -972891995;
assign addr[53437]= -904098143;
assign addr[53438]= -834157373;
assign addr[53439]= -763158411;
assign addr[53440]= -691191324;
assign addr[53441]= -618347408;
assign addr[53442]= -544719071;
assign addr[53443]= -470399716;
assign addr[53444]= -395483624;
assign addr[53445]= -320065829;
assign addr[53446]= -244242007;
assign addr[53447]= -168108346;
assign addr[53448]= -91761426;
assign addr[53449]= -15298099;
assign addr[53450]= 61184634;
assign addr[53451]= 137589750;
assign addr[53452]= 213820322;
assign addr[53453]= 289779648;
assign addr[53454]= 365371365;
assign addr[53455]= 440499581;
assign addr[53456]= 515068990;
assign addr[53457]= 588984994;
assign addr[53458]= 662153826;
assign addr[53459]= 734482665;
assign addr[53460]= 805879757;
assign addr[53461]= 876254528;
assign addr[53462]= 945517704;
assign addr[53463]= 1013581418;
assign addr[53464]= 1080359326;
assign addr[53465]= 1145766716;
assign addr[53466]= 1209720613;
assign addr[53467]= 1272139887;
assign addr[53468]= 1332945355;
assign addr[53469]= 1392059879;
assign addr[53470]= 1449408469;
assign addr[53471]= 1504918373;
assign addr[53472]= 1558519173;
assign addr[53473]= 1610142873;
assign addr[53474]= 1659723983;
assign addr[53475]= 1707199606;
assign addr[53476]= 1752509516;
assign addr[53477]= 1795596234;
assign addr[53478]= 1836405100;
assign addr[53479]= 1874884346;
assign addr[53480]= 1910985158;
assign addr[53481]= 1944661739;
assign addr[53482]= 1975871368;
assign addr[53483]= 2004574453;
assign addr[53484]= 2030734582;
assign addr[53485]= 2054318569;
assign addr[53486]= 2075296495;
assign addr[53487]= 2093641749;
assign addr[53488]= 2109331059;
assign addr[53489]= 2122344521;
assign addr[53490]= 2132665626;
assign addr[53491]= 2140281282;
assign addr[53492]= 2145181827;
assign addr[53493]= 2147361045;
assign addr[53494]= 2146816171;
assign addr[53495]= 2143547897;
assign addr[53496]= 2137560369;
assign addr[53497]= 2128861181;
assign addr[53498]= 2117461370;
assign addr[53499]= 2103375398;
assign addr[53500]= 2086621133;
assign addr[53501]= 2067219829;
assign addr[53502]= 2045196100;
assign addr[53503]= 2020577882;
assign addr[53504]= 1993396407;
assign addr[53505]= 1963686155;
assign addr[53506]= 1931484818;
assign addr[53507]= 1896833245;
assign addr[53508]= 1859775393;
assign addr[53509]= 1820358275;
assign addr[53510]= 1778631892;
assign addr[53511]= 1734649179;
assign addr[53512]= 1688465931;
assign addr[53513]= 1640140734;
assign addr[53514]= 1589734894;
assign addr[53515]= 1537312353;
assign addr[53516]= 1482939614;
assign addr[53517]= 1426685652;
assign addr[53518]= 1368621831;
assign addr[53519]= 1308821808;
assign addr[53520]= 1247361445;
assign addr[53521]= 1184318708;
assign addr[53522]= 1119773573;
assign addr[53523]= 1053807919;
assign addr[53524]= 986505429;
assign addr[53525]= 917951481;
assign addr[53526]= 848233042;
assign addr[53527]= 777438554;
assign addr[53528]= 705657826;
assign addr[53529]= 632981917;
assign addr[53530]= 559503022;
assign addr[53531]= 485314355;
assign addr[53532]= 410510029;
assign addr[53533]= 335184940;
assign addr[53534]= 259434643;
assign addr[53535]= 183355234;
assign addr[53536]= 107043224;
assign addr[53537]= 30595422;
assign addr[53538]= -45891193;
assign addr[53539]= -122319591;
assign addr[53540]= -198592817;
assign addr[53541]= -274614114;
assign addr[53542]= -350287041;
assign addr[53543]= -425515602;
assign addr[53544]= -500204365;
assign addr[53545]= -574258580;
assign addr[53546]= -647584304;
assign addr[53547]= -720088517;
assign addr[53548]= -791679244;
assign addr[53549]= -862265664;
assign addr[53550]= -931758235;
assign addr[53551]= -1000068799;
assign addr[53552]= -1067110699;
assign addr[53553]= -1132798888;
assign addr[53554]= -1197050035;
assign addr[53555]= -1259782632;
assign addr[53556]= -1320917099;
assign addr[53557]= -1380375881;
assign addr[53558]= -1438083551;
assign addr[53559]= -1493966902;
assign addr[53560]= -1547955041;
assign addr[53561]= -1599979481;
assign addr[53562]= -1649974225;
assign addr[53563]= -1697875851;
assign addr[53564]= -1743623590;
assign addr[53565]= -1787159411;
assign addr[53566]= -1828428082;
assign addr[53567]= -1867377253;
assign addr[53568]= -1903957513;
assign addr[53569]= -1938122457;
assign addr[53570]= -1969828744;
assign addr[53571]= -1999036154;
assign addr[53572]= -2025707632;
assign addr[53573]= -2049809346;
assign addr[53574]= -2071310720;
assign addr[53575]= -2090184478;
assign addr[53576]= -2106406677;
assign addr[53577]= -2119956737;
assign addr[53578]= -2130817471;
assign addr[53579]= -2138975100;
assign addr[53580]= -2144419275;
assign addr[53581]= -2147143090;
assign addr[53582]= -2147143090;
assign addr[53583]= -2144419275;
assign addr[53584]= -2138975100;
assign addr[53585]= -2130817471;
assign addr[53586]= -2119956737;
assign addr[53587]= -2106406677;
assign addr[53588]= -2090184478;
assign addr[53589]= -2071310720;
assign addr[53590]= -2049809346;
assign addr[53591]= -2025707632;
assign addr[53592]= -1999036154;
assign addr[53593]= -1969828744;
assign addr[53594]= -1938122457;
assign addr[53595]= -1903957513;
assign addr[53596]= -1867377253;
assign addr[53597]= -1828428082;
assign addr[53598]= -1787159411;
assign addr[53599]= -1743623590;
assign addr[53600]= -1697875851;
assign addr[53601]= -1649974225;
assign addr[53602]= -1599979481;
assign addr[53603]= -1547955041;
assign addr[53604]= -1493966902;
assign addr[53605]= -1438083551;
assign addr[53606]= -1380375881;
assign addr[53607]= -1320917099;
assign addr[53608]= -1259782632;
assign addr[53609]= -1197050035;
assign addr[53610]= -1132798888;
assign addr[53611]= -1067110699;
assign addr[53612]= -1000068799;
assign addr[53613]= -931758235;
assign addr[53614]= -862265664;
assign addr[53615]= -791679244;
assign addr[53616]= -720088517;
assign addr[53617]= -647584304;
assign addr[53618]= -574258580;
assign addr[53619]= -500204365;
assign addr[53620]= -425515602;
assign addr[53621]= -350287041;
assign addr[53622]= -274614114;
assign addr[53623]= -198592817;
assign addr[53624]= -122319591;
assign addr[53625]= -45891193;
assign addr[53626]= 30595422;
assign addr[53627]= 107043224;
assign addr[53628]= 183355234;
assign addr[53629]= 259434643;
assign addr[53630]= 335184940;
assign addr[53631]= 410510029;
assign addr[53632]= 485314355;
assign addr[53633]= 559503022;
assign addr[53634]= 632981917;
assign addr[53635]= 705657826;
assign addr[53636]= 777438554;
assign addr[53637]= 848233042;
assign addr[53638]= 917951481;
assign addr[53639]= 986505429;
assign addr[53640]= 1053807919;
assign addr[53641]= 1119773573;
assign addr[53642]= 1184318708;
assign addr[53643]= 1247361445;
assign addr[53644]= 1308821808;
assign addr[53645]= 1368621831;
assign addr[53646]= 1426685652;
assign addr[53647]= 1482939614;
assign addr[53648]= 1537312353;
assign addr[53649]= 1589734894;
assign addr[53650]= 1640140734;
assign addr[53651]= 1688465931;
assign addr[53652]= 1734649179;
assign addr[53653]= 1778631892;
assign addr[53654]= 1820358275;
assign addr[53655]= 1859775393;
assign addr[53656]= 1896833245;
assign addr[53657]= 1931484818;
assign addr[53658]= 1963686155;
assign addr[53659]= 1993396407;
assign addr[53660]= 2020577882;
assign addr[53661]= 2045196100;
assign addr[53662]= 2067219829;
assign addr[53663]= 2086621133;
assign addr[53664]= 2103375398;
assign addr[53665]= 2117461370;
assign addr[53666]= 2128861181;
assign addr[53667]= 2137560369;
assign addr[53668]= 2143547897;
assign addr[53669]= 2146816171;
assign addr[53670]= 2147361045;
assign addr[53671]= 2145181827;
assign addr[53672]= 2140281282;
assign addr[53673]= 2132665626;
assign addr[53674]= 2122344521;
assign addr[53675]= 2109331059;
assign addr[53676]= 2093641749;
assign addr[53677]= 2075296495;
assign addr[53678]= 2054318569;
assign addr[53679]= 2030734582;
assign addr[53680]= 2004574453;
assign addr[53681]= 1975871368;
assign addr[53682]= 1944661739;
assign addr[53683]= 1910985158;
assign addr[53684]= 1874884346;
assign addr[53685]= 1836405100;
assign addr[53686]= 1795596234;
assign addr[53687]= 1752509516;
assign addr[53688]= 1707199606;
assign addr[53689]= 1659723983;
assign addr[53690]= 1610142873;
assign addr[53691]= 1558519173;
assign addr[53692]= 1504918373;
assign addr[53693]= 1449408469;
assign addr[53694]= 1392059879;
assign addr[53695]= 1332945355;
assign addr[53696]= 1272139887;
assign addr[53697]= 1209720613;
assign addr[53698]= 1145766716;
assign addr[53699]= 1080359326;
assign addr[53700]= 1013581418;
assign addr[53701]= 945517704;
assign addr[53702]= 876254528;
assign addr[53703]= 805879757;
assign addr[53704]= 734482665;
assign addr[53705]= 662153826;
assign addr[53706]= 588984994;
assign addr[53707]= 515068990;
assign addr[53708]= 440499581;
assign addr[53709]= 365371365;
assign addr[53710]= 289779648;
assign addr[53711]= 213820322;
assign addr[53712]= 137589750;
assign addr[53713]= 61184634;
assign addr[53714]= -15298099;
assign addr[53715]= -91761426;
assign addr[53716]= -168108346;
assign addr[53717]= -244242007;
assign addr[53718]= -320065829;
assign addr[53719]= -395483624;
assign addr[53720]= -470399716;
assign addr[53721]= -544719071;
assign addr[53722]= -618347408;
assign addr[53723]= -691191324;
assign addr[53724]= -763158411;
assign addr[53725]= -834157373;
assign addr[53726]= -904098143;
assign addr[53727]= -972891995;
assign addr[53728]= -1040451659;
assign addr[53729]= -1106691431;
assign addr[53730]= -1171527280;
assign addr[53731]= -1234876957;
assign addr[53732]= -1296660098;
assign addr[53733]= -1356798326;
assign addr[53734]= -1415215352;
assign addr[53735]= -1471837070;
assign addr[53736]= -1526591649;
assign addr[53737]= -1579409630;
assign addr[53738]= -1630224009;
assign addr[53739]= -1678970324;
assign addr[53740]= -1725586737;
assign addr[53741]= -1770014111;
assign addr[53742]= -1812196087;
assign addr[53743]= -1852079154;
assign addr[53744]= -1889612716;
assign addr[53745]= -1924749160;
assign addr[53746]= -1957443913;
assign addr[53747]= -1987655498;
assign addr[53748]= -2015345591;
assign addr[53749]= -2040479063;
assign addr[53750]= -2063024031;
assign addr[53751]= -2082951896;
assign addr[53752]= -2100237377;
assign addr[53753]= -2114858546;
assign addr[53754]= -2126796855;
assign addr[53755]= -2136037160;
assign addr[53756]= -2142567738;
assign addr[53757]= -2146380306;
assign addr[53758]= -2147470025;
assign addr[53759]= -2145835515;
assign addr[53760]= -2141478848;
assign addr[53761]= -2134405552;
assign addr[53762]= -2124624598;
assign addr[53763]= -2112148396;
assign addr[53764]= -2096992772;
assign addr[53765]= -2079176953;
assign addr[53766]= -2058723538;
assign addr[53767]= -2035658475;
assign addr[53768]= -2010011024;
assign addr[53769]= -1981813720;
assign addr[53770]= -1951102334;
assign addr[53771]= -1917915825;
assign addr[53772]= -1882296293;
assign addr[53773]= -1844288924;
assign addr[53774]= -1803941934;
assign addr[53775]= -1761306505;
assign addr[53776]= -1716436725;
assign addr[53777]= -1669389513;
assign addr[53778]= -1620224553;
assign addr[53779]= -1569004214;
assign addr[53780]= -1515793473;
assign addr[53781]= -1460659832;
assign addr[53782]= -1403673233;
assign addr[53783]= -1344905966;
assign addr[53784]= -1284432584;
assign addr[53785]= -1222329801;
assign addr[53786]= -1158676398;
assign addr[53787]= -1093553126;
assign addr[53788]= -1027042599;
assign addr[53789]= -959229189;
assign addr[53790]= -890198924;
assign addr[53791]= -820039373;
assign addr[53792]= -748839539;
assign addr[53793]= -676689746;
assign addr[53794]= -603681519;
assign addr[53795]= -529907477;
assign addr[53796]= -455461206;
assign addr[53797]= -380437148;
assign addr[53798]= -304930476;
assign addr[53799]= -229036977;
assign addr[53800]= -152852926;
assign addr[53801]= -76474970;
assign addr[53802]= 0;
assign addr[53803]= 76474970;
assign addr[53804]= 152852926;
assign addr[53805]= 229036977;
assign addr[53806]= 304930476;
assign addr[53807]= 380437148;
assign addr[53808]= 455461206;
assign addr[53809]= 529907477;
assign addr[53810]= 603681519;
assign addr[53811]= 676689746;
assign addr[53812]= 748839539;
assign addr[53813]= 820039373;
assign addr[53814]= 890198924;
assign addr[53815]= 959229189;
assign addr[53816]= 1027042599;
assign addr[53817]= 1093553126;
assign addr[53818]= 1158676398;
assign addr[53819]= 1222329801;
assign addr[53820]= 1284432584;
assign addr[53821]= 1344905966;
assign addr[53822]= 1403673233;
assign addr[53823]= 1460659832;
assign addr[53824]= 1515793473;
assign addr[53825]= 1569004214;
assign addr[53826]= 1620224553;
assign addr[53827]= 1669389513;
assign addr[53828]= 1716436725;
assign addr[53829]= 1761306505;
assign addr[53830]= 1803941934;
assign addr[53831]= 1844288924;
assign addr[53832]= 1882296293;
assign addr[53833]= 1917915825;
assign addr[53834]= 1951102334;
assign addr[53835]= 1981813720;
assign addr[53836]= 2010011024;
assign addr[53837]= 2035658475;
assign addr[53838]= 2058723538;
assign addr[53839]= 2079176953;
assign addr[53840]= 2096992772;
assign addr[53841]= 2112148396;
assign addr[53842]= 2124624598;
assign addr[53843]= 2134405552;
assign addr[53844]= 2141478848;
assign addr[53845]= 2145835515;
assign addr[53846]= 2147470025;
assign addr[53847]= 2146380306;
assign addr[53848]= 2142567738;
assign addr[53849]= 2136037160;
assign addr[53850]= 2126796855;
assign addr[53851]= 2114858546;
assign addr[53852]= 2100237377;
assign addr[53853]= 2082951896;
assign addr[53854]= 2063024031;
assign addr[53855]= 2040479063;
assign addr[53856]= 2015345591;
assign addr[53857]= 1987655498;
assign addr[53858]= 1957443913;
assign addr[53859]= 1924749160;
assign addr[53860]= 1889612716;
assign addr[53861]= 1852079154;
assign addr[53862]= 1812196087;
assign addr[53863]= 1770014111;
assign addr[53864]= 1725586737;
assign addr[53865]= 1678970324;
assign addr[53866]= 1630224009;
assign addr[53867]= 1579409630;
assign addr[53868]= 1526591649;
assign addr[53869]= 1471837070;
assign addr[53870]= 1415215352;
assign addr[53871]= 1356798326;
assign addr[53872]= 1296660098;
assign addr[53873]= 1234876957;
assign addr[53874]= 1171527280;
assign addr[53875]= 1106691431;
assign addr[53876]= 1040451659;
assign addr[53877]= 972891995;
assign addr[53878]= 904098143;
assign addr[53879]= 834157373;
assign addr[53880]= 763158411;
assign addr[53881]= 691191324;
assign addr[53882]= 618347408;
assign addr[53883]= 544719071;
assign addr[53884]= 470399716;
assign addr[53885]= 395483624;
assign addr[53886]= 320065829;
assign addr[53887]= 244242007;
assign addr[53888]= 168108346;
assign addr[53889]= 91761426;
assign addr[53890]= 15298099;
assign addr[53891]= -61184634;
assign addr[53892]= -137589750;
assign addr[53893]= -213820322;
assign addr[53894]= -289779648;
assign addr[53895]= -365371365;
assign addr[53896]= -440499581;
assign addr[53897]= -515068990;
assign addr[53898]= -588984994;
assign addr[53899]= -662153826;
assign addr[53900]= -734482665;
assign addr[53901]= -805879757;
assign addr[53902]= -876254528;
assign addr[53903]= -945517704;
assign addr[53904]= -1013581418;
assign addr[53905]= -1080359326;
assign addr[53906]= -1145766716;
assign addr[53907]= -1209720613;
assign addr[53908]= -1272139887;
assign addr[53909]= -1332945355;
assign addr[53910]= -1392059879;
assign addr[53911]= -1449408469;
assign addr[53912]= -1504918373;
assign addr[53913]= -1558519173;
assign addr[53914]= -1610142873;
assign addr[53915]= -1659723983;
assign addr[53916]= -1707199606;
assign addr[53917]= -1752509516;
assign addr[53918]= -1795596234;
assign addr[53919]= -1836405100;
assign addr[53920]= -1874884346;
assign addr[53921]= -1910985158;
assign addr[53922]= -1944661739;
assign addr[53923]= -1975871368;
assign addr[53924]= -2004574453;
assign addr[53925]= -2030734582;
assign addr[53926]= -2054318569;
assign addr[53927]= -2075296495;
assign addr[53928]= -2093641749;
assign addr[53929]= -2109331059;
assign addr[53930]= -2122344521;
assign addr[53931]= -2132665626;
assign addr[53932]= -2140281282;
assign addr[53933]= -2145181827;
assign addr[53934]= -2147361045;
assign addr[53935]= -2146816171;
assign addr[53936]= -2143547897;
assign addr[53937]= -2137560369;
assign addr[53938]= -2128861181;
assign addr[53939]= -2117461370;
assign addr[53940]= -2103375398;
assign addr[53941]= -2086621133;
assign addr[53942]= -2067219829;
assign addr[53943]= -2045196100;
assign addr[53944]= -2020577882;
assign addr[53945]= -1993396407;
assign addr[53946]= -1963686155;
assign addr[53947]= -1931484818;
assign addr[53948]= -1896833245;
assign addr[53949]= -1859775393;
assign addr[53950]= -1820358275;
assign addr[53951]= -1778631892;
assign addr[53952]= -1734649179;
assign addr[53953]= -1688465931;
assign addr[53954]= -1640140734;
assign addr[53955]= -1589734894;
assign addr[53956]= -1537312353;
assign addr[53957]= -1482939614;
assign addr[53958]= -1426685652;
assign addr[53959]= -1368621831;
assign addr[53960]= -1308821808;
assign addr[53961]= -1247361445;
assign addr[53962]= -1184318708;
assign addr[53963]= -1119773573;
assign addr[53964]= -1053807919;
assign addr[53965]= -986505429;
assign addr[53966]= -917951481;
assign addr[53967]= -848233042;
assign addr[53968]= -777438554;
assign addr[53969]= -705657826;
assign addr[53970]= -632981917;
assign addr[53971]= -559503022;
assign addr[53972]= -485314355;
assign addr[53973]= -410510029;
assign addr[53974]= -335184940;
assign addr[53975]= -259434643;
assign addr[53976]= -183355234;
assign addr[53977]= -107043224;
assign addr[53978]= -30595422;
assign addr[53979]= 45891193;
assign addr[53980]= 122319591;
assign addr[53981]= 198592817;
assign addr[53982]= 274614114;
assign addr[53983]= 350287041;
assign addr[53984]= 425515602;
assign addr[53985]= 500204365;
assign addr[53986]= 574258580;
assign addr[53987]= 647584304;
assign addr[53988]= 720088517;
assign addr[53989]= 791679244;
assign addr[53990]= 862265664;
assign addr[53991]= 931758235;
assign addr[53992]= 1000068799;
assign addr[53993]= 1067110699;
assign addr[53994]= 1132798888;
assign addr[53995]= 1197050035;
assign addr[53996]= 1259782632;
assign addr[53997]= 1320917099;
assign addr[53998]= 1380375881;
assign addr[53999]= 1438083551;
assign addr[54000]= 1493966902;
assign addr[54001]= 1547955041;
assign addr[54002]= 1599979481;
assign addr[54003]= 1649974225;
assign addr[54004]= 1697875851;
assign addr[54005]= 1743623590;
assign addr[54006]= 1787159411;
assign addr[54007]= 1828428082;
assign addr[54008]= 1867377253;
assign addr[54009]= 1903957513;
assign addr[54010]= 1938122457;
assign addr[54011]= 1969828744;
assign addr[54012]= 1999036154;
assign addr[54013]= 2025707632;
assign addr[54014]= 2049809346;
assign addr[54015]= 2071310720;
assign addr[54016]= 2090184478;
assign addr[54017]= 2106406677;
assign addr[54018]= 2119956737;
assign addr[54019]= 2130817471;
assign addr[54020]= 2138975100;
assign addr[54021]= 2144419275;
assign addr[54022]= 2147143090;
assign addr[54023]= 2147143090;
assign addr[54024]= 2144419275;
assign addr[54025]= 2138975100;
assign addr[54026]= 2130817471;
assign addr[54027]= 2119956737;
assign addr[54028]= 2106406677;
assign addr[54029]= 2090184478;
assign addr[54030]= 2071310720;
assign addr[54031]= 2049809346;
assign addr[54032]= 2025707632;
assign addr[54033]= 1999036154;
assign addr[54034]= 1969828744;
assign addr[54035]= 1938122457;
assign addr[54036]= 1903957513;
assign addr[54037]= 1867377253;
assign addr[54038]= 1828428082;
assign addr[54039]= 1787159411;
assign addr[54040]= 1743623590;
assign addr[54041]= 1697875851;
assign addr[54042]= 1649974225;
assign addr[54043]= 1599979481;
assign addr[54044]= 1547955041;
assign addr[54045]= 1493966902;
assign addr[54046]= 1438083551;
assign addr[54047]= 1380375881;
assign addr[54048]= 1320917099;
assign addr[54049]= 1259782632;
assign addr[54050]= 1197050035;
assign addr[54051]= 1132798888;
assign addr[54052]= 1067110699;
assign addr[54053]= 1000068799;
assign addr[54054]= 931758235;
assign addr[54055]= 862265664;
assign addr[54056]= 791679244;
assign addr[54057]= 720088517;
assign addr[54058]= 647584304;
assign addr[54059]= 574258580;
assign addr[54060]= 500204365;
assign addr[54061]= 425515602;
assign addr[54062]= 350287041;
assign addr[54063]= 274614114;
assign addr[54064]= 198592817;
assign addr[54065]= 122319591;
assign addr[54066]= 45891193;
assign addr[54067]= -30595422;
assign addr[54068]= -107043224;
assign addr[54069]= -183355234;
assign addr[54070]= -259434643;
assign addr[54071]= -335184940;
assign addr[54072]= -410510029;
assign addr[54073]= -485314355;
assign addr[54074]= -559503022;
assign addr[54075]= -632981917;
assign addr[54076]= -705657826;
assign addr[54077]= -777438554;
assign addr[54078]= -848233042;
assign addr[54079]= -917951481;
assign addr[54080]= -986505429;
assign addr[54081]= -1053807919;
assign addr[54082]= -1119773573;
assign addr[54083]= -1184318708;
assign addr[54084]= -1247361445;
assign addr[54085]= -1308821808;
assign addr[54086]= -1368621831;
assign addr[54087]= -1426685652;
assign addr[54088]= -1482939614;
assign addr[54089]= -1537312353;
assign addr[54090]= -1589734894;
assign addr[54091]= -1640140734;
assign addr[54092]= -1688465931;
assign addr[54093]= -1734649179;
assign addr[54094]= -1778631892;
assign addr[54095]= -1820358275;
assign addr[54096]= -1859775393;
assign addr[54097]= -1896833245;
assign addr[54098]= -1931484818;
assign addr[54099]= -1963686155;
assign addr[54100]= -1993396407;
assign addr[54101]= -2020577882;
assign addr[54102]= -2045196100;
assign addr[54103]= -2067219829;
assign addr[54104]= -2086621133;
assign addr[54105]= -2103375398;
assign addr[54106]= -2117461370;
assign addr[54107]= -2128861181;
assign addr[54108]= -2137560369;
assign addr[54109]= -2143547897;
assign addr[54110]= -2146816171;
assign addr[54111]= -2147361045;
assign addr[54112]= -2145181827;
assign addr[54113]= -2140281282;
assign addr[54114]= -2132665626;
assign addr[54115]= -2122344521;
assign addr[54116]= -2109331059;
assign addr[54117]= -2093641749;
assign addr[54118]= -2075296495;
assign addr[54119]= -2054318569;
assign addr[54120]= -2030734582;
assign addr[54121]= -2004574453;
assign addr[54122]= -1975871368;
assign addr[54123]= -1944661739;
assign addr[54124]= -1910985158;
assign addr[54125]= -1874884346;
assign addr[54126]= -1836405100;
assign addr[54127]= -1795596234;
assign addr[54128]= -1752509516;
assign addr[54129]= -1707199606;
assign addr[54130]= -1659723983;
assign addr[54131]= -1610142873;
assign addr[54132]= -1558519173;
assign addr[54133]= -1504918373;
assign addr[54134]= -1449408469;
assign addr[54135]= -1392059879;
assign addr[54136]= -1332945355;
assign addr[54137]= -1272139887;
assign addr[54138]= -1209720613;
assign addr[54139]= -1145766716;
assign addr[54140]= -1080359326;
assign addr[54141]= -1013581418;
assign addr[54142]= -945517704;
assign addr[54143]= -876254528;
assign addr[54144]= -805879757;
assign addr[54145]= -734482665;
assign addr[54146]= -662153826;
assign addr[54147]= -588984994;
assign addr[54148]= -515068990;
assign addr[54149]= -440499581;
assign addr[54150]= -365371365;
assign addr[54151]= -289779648;
assign addr[54152]= -213820322;
assign addr[54153]= -137589750;
assign addr[54154]= -61184634;
assign addr[54155]= 15298099;
assign addr[54156]= 91761426;
assign addr[54157]= 168108346;
assign addr[54158]= 244242007;
assign addr[54159]= 320065829;
assign addr[54160]= 395483624;
assign addr[54161]= 470399716;
assign addr[54162]= 544719071;
assign addr[54163]= 618347408;
assign addr[54164]= 691191324;
assign addr[54165]= 763158411;
assign addr[54166]= 834157373;
assign addr[54167]= 904098143;
assign addr[54168]= 972891995;
assign addr[54169]= 1040451659;
assign addr[54170]= 1106691431;
assign addr[54171]= 1171527280;
assign addr[54172]= 1234876957;
assign addr[54173]= 1296660098;
assign addr[54174]= 1356798326;
assign addr[54175]= 1415215352;
assign addr[54176]= 1471837070;
assign addr[54177]= 1526591649;
assign addr[54178]= 1579409630;
assign addr[54179]= 1630224009;
assign addr[54180]= 1678970324;
assign addr[54181]= 1725586737;
assign addr[54182]= 1770014111;
assign addr[54183]= 1812196087;
assign addr[54184]= 1852079154;
assign addr[54185]= 1889612716;
assign addr[54186]= 1924749160;
assign addr[54187]= 1957443913;
assign addr[54188]= 1987655498;
assign addr[54189]= 2015345591;
assign addr[54190]= 2040479063;
assign addr[54191]= 2063024031;
assign addr[54192]= 2082951896;
assign addr[54193]= 2100237377;
assign addr[54194]= 2114858546;
assign addr[54195]= 2126796855;
assign addr[54196]= 2136037160;
assign addr[54197]= 2142567738;
assign addr[54198]= 2146380306;
assign addr[54199]= 2147470025;
assign addr[54200]= 2145835515;
assign addr[54201]= 2141478848;
assign addr[54202]= 2134405552;
assign addr[54203]= 2124624598;
assign addr[54204]= 2112148396;
assign addr[54205]= 2096992772;
assign addr[54206]= 2079176953;
assign addr[54207]= 2058723538;
assign addr[54208]= 2035658475;
assign addr[54209]= 2010011024;
assign addr[54210]= 1981813720;
assign addr[54211]= 1951102334;
assign addr[54212]= 1917915825;
assign addr[54213]= 1882296293;
assign addr[54214]= 1844288924;
assign addr[54215]= 1803941934;
assign addr[54216]= 1761306505;
assign addr[54217]= 1716436725;
assign addr[54218]= 1669389513;
assign addr[54219]= 1620224553;
assign addr[54220]= 1569004214;
assign addr[54221]= 1515793473;
assign addr[54222]= 1460659832;
assign addr[54223]= 1403673233;
assign addr[54224]= 1344905966;
assign addr[54225]= 1284432584;
assign addr[54226]= 1222329801;
assign addr[54227]= 1158676398;
assign addr[54228]= 1093553126;
assign addr[54229]= 1027042599;
assign addr[54230]= 959229189;
assign addr[54231]= 890198924;
assign addr[54232]= 820039373;
assign addr[54233]= 748839539;
assign addr[54234]= 676689746;
assign addr[54235]= 603681519;
assign addr[54236]= 529907477;
assign addr[54237]= 455461206;
assign addr[54238]= 380437148;
assign addr[54239]= 304930476;
assign addr[54240]= 229036977;
assign addr[54241]= 152852926;
assign addr[54242]= 76474970;
assign addr[54243]= 0;
assign addr[54244]= -76474970;
assign addr[54245]= -152852926;
assign addr[54246]= -229036977;
assign addr[54247]= -304930476;
assign addr[54248]= -380437148;
assign addr[54249]= -455461206;
assign addr[54250]= -529907477;
assign addr[54251]= -603681519;
assign addr[54252]= -676689746;
assign addr[54253]= -748839539;
assign addr[54254]= -820039373;
assign addr[54255]= -890198924;
assign addr[54256]= -959229189;
assign addr[54257]= -1027042599;
assign addr[54258]= -1093553126;
assign addr[54259]= -1158676398;
assign addr[54260]= -1222329801;
assign addr[54261]= -1284432584;
assign addr[54262]= -1344905966;
assign addr[54263]= -1403673233;
assign addr[54264]= -1460659832;
assign addr[54265]= -1515793473;
assign addr[54266]= -1569004214;
assign addr[54267]= -1620224553;
assign addr[54268]= -1669389513;
assign addr[54269]= -1716436725;
assign addr[54270]= -1761306505;
assign addr[54271]= -1803941934;
assign addr[54272]= -1844288924;
assign addr[54273]= -1882296293;
assign addr[54274]= -1917915825;
assign addr[54275]= -1951102334;
assign addr[54276]= -1981813720;
assign addr[54277]= -2010011024;
assign addr[54278]= -2035658475;
assign addr[54279]= -2058723538;
assign addr[54280]= -2079176953;
assign addr[54281]= -2096992772;
assign addr[54282]= -2112148396;
assign addr[54283]= -2124624598;
assign addr[54284]= -2134405552;
assign addr[54285]= -2141478848;
assign addr[54286]= -2145835515;
assign addr[54287]= -2147470025;
assign addr[54288]= -2146380306;
assign addr[54289]= -2142567738;
assign addr[54290]= -2136037160;
assign addr[54291]= -2126796855;
assign addr[54292]= -2114858546;
assign addr[54293]= -2100237377;
assign addr[54294]= -2082951896;
assign addr[54295]= -2063024031;
assign addr[54296]= -2040479063;
assign addr[54297]= -2015345591;
assign addr[54298]= -1987655498;
assign addr[54299]= -1957443913;
assign addr[54300]= -1924749160;
assign addr[54301]= -1889612716;
assign addr[54302]= -1852079154;
assign addr[54303]= -1812196087;
assign addr[54304]= -1770014111;
assign addr[54305]= -1725586737;
assign addr[54306]= -1678970324;
assign addr[54307]= -1630224009;
assign addr[54308]= -1579409630;
assign addr[54309]= -1526591649;
assign addr[54310]= -1471837070;
assign addr[54311]= -1415215352;
assign addr[54312]= -1356798326;
assign addr[54313]= -1296660098;
assign addr[54314]= -1234876957;
assign addr[54315]= -1171527280;
assign addr[54316]= -1106691431;
assign addr[54317]= -1040451659;
assign addr[54318]= -972891995;
assign addr[54319]= -904098143;
assign addr[54320]= -834157373;
assign addr[54321]= -763158411;
assign addr[54322]= -691191324;
assign addr[54323]= -618347408;
assign addr[54324]= -544719071;
assign addr[54325]= -470399716;
assign addr[54326]= -395483624;
assign addr[54327]= -320065829;
assign addr[54328]= -244242007;
assign addr[54329]= -168108346;
assign addr[54330]= -91761426;
assign addr[54331]= -15298099;
assign addr[54332]= 61184634;
assign addr[54333]= 137589750;
assign addr[54334]= 213820322;
assign addr[54335]= 289779648;
assign addr[54336]= 365371365;
assign addr[54337]= 440499581;
assign addr[54338]= 515068990;
assign addr[54339]= 588984994;
assign addr[54340]= 662153826;
assign addr[54341]= 734482665;
assign addr[54342]= 805879757;
assign addr[54343]= 876254528;
assign addr[54344]= 945517704;
assign addr[54345]= 1013581418;
assign addr[54346]= 1080359326;
assign addr[54347]= 1145766716;
assign addr[54348]= 1209720613;
assign addr[54349]= 1272139887;
assign addr[54350]= 1332945355;
assign addr[54351]= 1392059879;
assign addr[54352]= 1449408469;
assign addr[54353]= 1504918373;
assign addr[54354]= 1558519173;
assign addr[54355]= 1610142873;
assign addr[54356]= 1659723983;
assign addr[54357]= 1707199606;
assign addr[54358]= 1752509516;
assign addr[54359]= 1795596234;
assign addr[54360]= 1836405100;
assign addr[54361]= 1874884346;
assign addr[54362]= 1910985158;
assign addr[54363]= 1944661739;
assign addr[54364]= 1975871368;
assign addr[54365]= 2004574453;
assign addr[54366]= 2030734582;
assign addr[54367]= 2054318569;
assign addr[54368]= 2075296495;
assign addr[54369]= 2093641749;
assign addr[54370]= 2109331059;
assign addr[54371]= 2122344521;
assign addr[54372]= 2132665626;
assign addr[54373]= 2140281282;
assign addr[54374]= 2145181827;
assign addr[54375]= 2147361045;
assign addr[54376]= 2146816171;
assign addr[54377]= 2143547897;
assign addr[54378]= 2137560369;
assign addr[54379]= 2128861181;
assign addr[54380]= 2117461370;
assign addr[54381]= 2103375398;
assign addr[54382]= 2086621133;
assign addr[54383]= 2067219829;
assign addr[54384]= 2045196100;
assign addr[54385]= 2020577882;
assign addr[54386]= 1993396407;
assign addr[54387]= 1963686155;
assign addr[54388]= 1931484818;
assign addr[54389]= 1896833245;
assign addr[54390]= 1859775393;
assign addr[54391]= 1820358275;
assign addr[54392]= 1778631892;
assign addr[54393]= 1734649179;
assign addr[54394]= 1688465931;
assign addr[54395]= 1640140734;
assign addr[54396]= 1589734894;
assign addr[54397]= 1537312353;
assign addr[54398]= 1482939614;
assign addr[54399]= 1426685652;
assign addr[54400]= 1368621831;
assign addr[54401]= 1308821808;
assign addr[54402]= 1247361445;
assign addr[54403]= 1184318708;
assign addr[54404]= 1119773573;
assign addr[54405]= 1053807919;
assign addr[54406]= 986505429;
assign addr[54407]= 917951481;
assign addr[54408]= 848233042;
assign addr[54409]= 777438554;
assign addr[54410]= 705657826;
assign addr[54411]= 632981917;
assign addr[54412]= 559503022;
assign addr[54413]= 485314355;
assign addr[54414]= 410510029;
assign addr[54415]= 335184940;
assign addr[54416]= 259434643;
assign addr[54417]= 183355234;
assign addr[54418]= 107043224;
assign addr[54419]= 30595422;
assign addr[54420]= -45891193;
assign addr[54421]= -122319591;
assign addr[54422]= -198592817;
assign addr[54423]= -274614114;
assign addr[54424]= -350287041;
assign addr[54425]= -425515602;
assign addr[54426]= -500204365;
assign addr[54427]= -574258580;
assign addr[54428]= -647584304;
assign addr[54429]= -720088517;
assign addr[54430]= -791679244;
assign addr[54431]= -862265664;
assign addr[54432]= -931758235;
assign addr[54433]= -1000068799;
assign addr[54434]= -1067110699;
assign addr[54435]= -1132798888;
assign addr[54436]= -1197050035;
assign addr[54437]= -1259782632;
assign addr[54438]= -1320917099;
assign addr[54439]= -1380375881;
assign addr[54440]= -1438083551;
assign addr[54441]= -1493966902;
assign addr[54442]= -1547955041;
assign addr[54443]= -1599979481;
assign addr[54444]= -1649974225;
assign addr[54445]= -1697875851;
assign addr[54446]= -1743623590;
assign addr[54447]= -1787159411;
assign addr[54448]= -1828428082;
assign addr[54449]= -1867377253;
assign addr[54450]= -1903957513;
assign addr[54451]= -1938122457;
assign addr[54452]= -1969828744;
assign addr[54453]= -1999036154;
assign addr[54454]= -2025707632;
assign addr[54455]= -2049809346;
assign addr[54456]= -2071310720;
assign addr[54457]= -2090184478;
assign addr[54458]= -2106406677;
assign addr[54459]= -2119956737;
assign addr[54460]= -2130817471;
assign addr[54461]= -2138975100;
assign addr[54462]= -2144419275;
assign addr[54463]= -2147143090;
assign addr[54464]= -2147143090;
assign addr[54465]= -2144419275;
assign addr[54466]= -2138975100;
assign addr[54467]= -2130817471;
assign addr[54468]= -2119956737;
assign addr[54469]= -2106406677;
assign addr[54470]= -2090184478;
assign addr[54471]= -2071310720;
assign addr[54472]= -2049809346;
assign addr[54473]= -2025707632;
assign addr[54474]= -1999036154;
assign addr[54475]= -1969828744;
assign addr[54476]= -1938122457;
assign addr[54477]= -1903957513;
assign addr[54478]= -1867377253;
assign addr[54479]= -1828428082;
assign addr[54480]= -1787159411;
assign addr[54481]= -1743623590;
assign addr[54482]= -1697875851;
assign addr[54483]= -1649974225;
assign addr[54484]= -1599979481;
assign addr[54485]= -1547955041;
assign addr[54486]= -1493966902;
assign addr[54487]= -1438083551;
assign addr[54488]= -1380375881;
assign addr[54489]= -1320917099;
assign addr[54490]= -1259782632;
assign addr[54491]= -1197050035;
assign addr[54492]= -1132798888;
assign addr[54493]= -1067110699;
assign addr[54494]= -1000068799;
assign addr[54495]= -931758235;
assign addr[54496]= -862265664;
assign addr[54497]= -791679244;
assign addr[54498]= -720088517;
assign addr[54499]= -647584304;
assign addr[54500]= -574258580;
assign addr[54501]= -500204365;
assign addr[54502]= -425515602;
assign addr[54503]= -350287041;
assign addr[54504]= -274614114;
assign addr[54505]= -198592817;
assign addr[54506]= -122319591;
assign addr[54507]= -45891193;
assign addr[54508]= 30595422;
assign addr[54509]= 107043224;
assign addr[54510]= 183355234;
assign addr[54511]= 259434643;
assign addr[54512]= 335184940;
assign addr[54513]= 410510029;
assign addr[54514]= 485314355;
assign addr[54515]= 559503022;
assign addr[54516]= 632981917;
assign addr[54517]= 705657826;
assign addr[54518]= 777438554;
assign addr[54519]= 848233042;
assign addr[54520]= 917951481;
assign addr[54521]= 986505429;
assign addr[54522]= 1053807919;
assign addr[54523]= 1119773573;
assign addr[54524]= 1184318708;
assign addr[54525]= 1247361445;
assign addr[54526]= 1308821808;
assign addr[54527]= 1368621831;
assign addr[54528]= 1426685652;
assign addr[54529]= 1482939614;
assign addr[54530]= 1537312353;
assign addr[54531]= 1589734894;
assign addr[54532]= 1640140734;
assign addr[54533]= 1688465931;
assign addr[54534]= 1734649179;
assign addr[54535]= 1778631892;
assign addr[54536]= 1820358275;
assign addr[54537]= 1859775393;
assign addr[54538]= 1896833245;
assign addr[54539]= 1931484818;
assign addr[54540]= 1963686155;
assign addr[54541]= 1993396407;
assign addr[54542]= 2020577882;
assign addr[54543]= 2045196100;
assign addr[54544]= 2067219829;
assign addr[54545]= 2086621133;
assign addr[54546]= 2103375398;
assign addr[54547]= 2117461370;
assign addr[54548]= 2128861181;
assign addr[54549]= 2137560369;
assign addr[54550]= 2143547897;
assign addr[54551]= 2146816171;
assign addr[54552]= 2147361045;
assign addr[54553]= 2145181827;
assign addr[54554]= 2140281282;
assign addr[54555]= 2132665626;
assign addr[54556]= 2122344521;
assign addr[54557]= 2109331059;
assign addr[54558]= 2093641749;
assign addr[54559]= 2075296495;
assign addr[54560]= 2054318569;
assign addr[54561]= 2030734582;
assign addr[54562]= 2004574453;
assign addr[54563]= 1975871368;
assign addr[54564]= 1944661739;
assign addr[54565]= 1910985158;
assign addr[54566]= 1874884346;
assign addr[54567]= 1836405100;
assign addr[54568]= 1795596234;
assign addr[54569]= 1752509516;
assign addr[54570]= 1707199606;
assign addr[54571]= 1659723983;
assign addr[54572]= 1610142873;
assign addr[54573]= 1558519173;
assign addr[54574]= 1504918373;
assign addr[54575]= 1449408469;
assign addr[54576]= 1392059879;
assign addr[54577]= 1332945355;
assign addr[54578]= 1272139887;
assign addr[54579]= 1209720613;
assign addr[54580]= 1145766716;
assign addr[54581]= 1080359326;
assign addr[54582]= 1013581418;
assign addr[54583]= 945517704;
assign addr[54584]= 876254528;
assign addr[54585]= 805879757;
assign addr[54586]= 734482665;
assign addr[54587]= 662153826;
assign addr[54588]= 588984994;
assign addr[54589]= 515068990;
assign addr[54590]= 440499581;
assign addr[54591]= 365371365;
assign addr[54592]= 289779648;
assign addr[54593]= 213820322;
assign addr[54594]= 137589750;
assign addr[54595]= 61184634;
assign addr[54596]= -15298099;
assign addr[54597]= -91761426;
assign addr[54598]= -168108346;
assign addr[54599]= -244242007;
assign addr[54600]= -320065829;
assign addr[54601]= -395483624;
assign addr[54602]= -470399716;
assign addr[54603]= -544719071;
assign addr[54604]= -618347408;
assign addr[54605]= -691191324;
assign addr[54606]= -763158411;
assign addr[54607]= -834157373;
assign addr[54608]= -904098143;
assign addr[54609]= -972891995;
assign addr[54610]= -1040451659;
assign addr[54611]= -1106691431;
assign addr[54612]= -1171527280;
assign addr[54613]= -1234876957;
assign addr[54614]= -1296660098;
assign addr[54615]= -1356798326;
assign addr[54616]= -1415215352;
assign addr[54617]= -1471837070;
assign addr[54618]= -1526591649;
assign addr[54619]= -1579409630;
assign addr[54620]= -1630224009;
assign addr[54621]= -1678970324;
assign addr[54622]= -1725586737;
assign addr[54623]= -1770014111;
assign addr[54624]= -1812196087;
assign addr[54625]= -1852079154;
assign addr[54626]= -1889612716;
assign addr[54627]= -1924749160;
assign addr[54628]= -1957443913;
assign addr[54629]= -1987655498;
assign addr[54630]= -2015345591;
assign addr[54631]= -2040479063;
assign addr[54632]= -2063024031;
assign addr[54633]= -2082951896;
assign addr[54634]= -2100237377;
assign addr[54635]= -2114858546;
assign addr[54636]= -2126796855;
assign addr[54637]= -2136037160;
assign addr[54638]= -2142567738;
assign addr[54639]= -2146380306;
assign addr[54640]= -2147470025;
assign addr[54641]= -2145835515;
assign addr[54642]= -2141478848;
assign addr[54643]= -2134405552;
assign addr[54644]= -2124624598;
assign addr[54645]= -2112148396;
assign addr[54646]= -2096992772;
assign addr[54647]= -2079176953;
assign addr[54648]= -2058723538;
assign addr[54649]= -2035658475;
assign addr[54650]= -2010011024;
assign addr[54651]= -1981813720;
assign addr[54652]= -1951102334;
assign addr[54653]= -1917915825;
assign addr[54654]= -1882296293;
assign addr[54655]= -1844288924;
assign addr[54656]= -1803941934;
assign addr[54657]= -1761306505;
assign addr[54658]= -1716436725;
assign addr[54659]= -1669389513;
assign addr[54660]= -1620224553;
assign addr[54661]= -1569004214;
assign addr[54662]= -1515793473;
assign addr[54663]= -1460659832;
assign addr[54664]= -1403673233;
assign addr[54665]= -1344905966;
assign addr[54666]= -1284432584;
assign addr[54667]= -1222329801;
assign addr[54668]= -1158676398;
assign addr[54669]= -1093553126;
assign addr[54670]= -1027042599;
assign addr[54671]= -959229189;
assign addr[54672]= -890198924;
assign addr[54673]= -820039373;
assign addr[54674]= -748839539;
assign addr[54675]= -676689746;
assign addr[54676]= -603681519;
assign addr[54677]= -529907477;
assign addr[54678]= -455461206;
assign addr[54679]= -380437148;
assign addr[54680]= -304930476;
assign addr[54681]= -229036977;
assign addr[54682]= -152852926;
assign addr[54683]= -76474970;
assign addr[54684]= 0;
assign addr[54685]= 76474970;
assign addr[54686]= 152852926;
assign addr[54687]= 229036977;
assign addr[54688]= 304930476;
assign addr[54689]= 380437148;
assign addr[54690]= 455461206;
assign addr[54691]= 529907477;
assign addr[54692]= 603681519;
assign addr[54693]= 676689746;
assign addr[54694]= 748839539;
assign addr[54695]= 820039373;
assign addr[54696]= 890198924;
assign addr[54697]= 959229189;
assign addr[54698]= 1027042599;
assign addr[54699]= 1093553126;
assign addr[54700]= 1158676398;
assign addr[54701]= 1222329801;
assign addr[54702]= 1284432584;
assign addr[54703]= 1344905966;
assign addr[54704]= 1403673233;
assign addr[54705]= 1460659832;
assign addr[54706]= 1515793473;
assign addr[54707]= 1569004214;
assign addr[54708]= 1620224553;
assign addr[54709]= 1669389513;
assign addr[54710]= 1716436725;
assign addr[54711]= 1761306505;
assign addr[54712]= 1803941934;
assign addr[54713]= 1844288924;
assign addr[54714]= 1882296293;
assign addr[54715]= 1917915825;
assign addr[54716]= 1951102334;
assign addr[54717]= 1981813720;
assign addr[54718]= 2010011024;
assign addr[54719]= 2035658475;
assign addr[54720]= 2058723538;
assign addr[54721]= 2079176953;
assign addr[54722]= 2096992772;
assign addr[54723]= 2112148396;
assign addr[54724]= 2124624598;
assign addr[54725]= 2134405552;
assign addr[54726]= 2141478848;
assign addr[54727]= 2145835515;
assign addr[54728]= 2147470025;
assign addr[54729]= 2146380306;
assign addr[54730]= 2142567738;
assign addr[54731]= 2136037160;
assign addr[54732]= 2126796855;
assign addr[54733]= 2114858546;
assign addr[54734]= 2100237377;
assign addr[54735]= 2082951896;
assign addr[54736]= 2063024031;
assign addr[54737]= 2040479063;
assign addr[54738]= 2015345591;
assign addr[54739]= 1987655498;
assign addr[54740]= 1957443913;
assign addr[54741]= 1924749160;
assign addr[54742]= 1889612716;
assign addr[54743]= 1852079154;
assign addr[54744]= 1812196087;
assign addr[54745]= 1770014111;
assign addr[54746]= 1725586737;
assign addr[54747]= 1678970324;
assign addr[54748]= 1630224009;
assign addr[54749]= 1579409630;
assign addr[54750]= 1526591649;
assign addr[54751]= 1471837070;
assign addr[54752]= 1415215352;
assign addr[54753]= 1356798326;
assign addr[54754]= 1296660098;
assign addr[54755]= 1234876957;
assign addr[54756]= 1171527280;
assign addr[54757]= 1106691431;
assign addr[54758]= 1040451659;
assign addr[54759]= 972891995;
assign addr[54760]= 904098143;
assign addr[54761]= 834157373;
assign addr[54762]= 763158411;
assign addr[54763]= 691191324;
assign addr[54764]= 618347408;
assign addr[54765]= 544719071;
assign addr[54766]= 470399716;
assign addr[54767]= 395483624;
assign addr[54768]= 320065829;
assign addr[54769]= 244242007;
assign addr[54770]= 168108346;
assign addr[54771]= 91761426;
assign addr[54772]= 15298099;
assign addr[54773]= -61184634;
assign addr[54774]= -137589750;
assign addr[54775]= -213820322;
assign addr[54776]= -289779648;
assign addr[54777]= -365371365;
assign addr[54778]= -440499581;
assign addr[54779]= -515068990;
assign addr[54780]= -588984994;
assign addr[54781]= -662153826;
assign addr[54782]= -734482665;
assign addr[54783]= -805879757;
assign addr[54784]= -876254528;
assign addr[54785]= -945517704;
assign addr[54786]= -1013581418;
assign addr[54787]= -1080359326;
assign addr[54788]= -1145766716;
assign addr[54789]= -1209720613;
assign addr[54790]= -1272139887;
assign addr[54791]= -1332945355;
assign addr[54792]= -1392059879;
assign addr[54793]= -1449408469;
assign addr[54794]= -1504918373;
assign addr[54795]= -1558519173;
assign addr[54796]= -1610142873;
assign addr[54797]= -1659723983;
assign addr[54798]= -1707199606;
assign addr[54799]= -1752509516;
assign addr[54800]= -1795596234;
assign addr[54801]= -1836405100;
assign addr[54802]= -1874884346;
assign addr[54803]= -1910985158;
assign addr[54804]= -1944661739;
assign addr[54805]= -1975871368;
assign addr[54806]= -2004574453;
assign addr[54807]= -2030734582;
assign addr[54808]= -2054318569;
assign addr[54809]= -2075296495;
assign addr[54810]= -2093641749;
assign addr[54811]= -2109331059;
assign addr[54812]= -2122344521;
assign addr[54813]= -2132665626;
assign addr[54814]= -2140281282;
assign addr[54815]= -2145181827;
assign addr[54816]= -2147361045;
assign addr[54817]= -2146816171;
assign addr[54818]= -2143547897;
assign addr[54819]= -2137560369;
assign addr[54820]= -2128861181;
assign addr[54821]= -2117461370;
assign addr[54822]= -2103375398;
assign addr[54823]= -2086621133;
assign addr[54824]= -2067219829;
assign addr[54825]= -2045196100;
assign addr[54826]= -2020577882;
assign addr[54827]= -1993396407;
assign addr[54828]= -1963686155;
assign addr[54829]= -1931484818;
assign addr[54830]= -1896833245;
assign addr[54831]= -1859775393;
assign addr[54832]= -1820358275;
assign addr[54833]= -1778631892;
assign addr[54834]= -1734649179;
assign addr[54835]= -1688465931;
assign addr[54836]= -1640140734;
assign addr[54837]= -1589734894;
assign addr[54838]= -1537312353;
assign addr[54839]= -1482939614;
assign addr[54840]= -1426685652;
assign addr[54841]= -1368621831;
assign addr[54842]= -1308821808;
assign addr[54843]= -1247361445;
assign addr[54844]= -1184318708;
assign addr[54845]= -1119773573;
assign addr[54846]= -1053807919;
assign addr[54847]= -986505429;
assign addr[54848]= -917951481;
assign addr[54849]= -848233042;
assign addr[54850]= -777438554;
assign addr[54851]= -705657826;
assign addr[54852]= -632981917;
assign addr[54853]= -559503022;
assign addr[54854]= -485314355;
assign addr[54855]= -410510029;
assign addr[54856]= -335184940;
assign addr[54857]= -259434643;
assign addr[54858]= -183355234;
assign addr[54859]= -107043224;
assign addr[54860]= -30595422;
assign addr[54861]= 45891193;
assign addr[54862]= 122319591;
assign addr[54863]= 198592817;
assign addr[54864]= 274614114;
assign addr[54865]= 350287041;
assign addr[54866]= 425515602;
assign addr[54867]= 500204365;
assign addr[54868]= 574258580;
assign addr[54869]= 647584304;
assign addr[54870]= 720088517;
assign addr[54871]= 791679244;
assign addr[54872]= 862265664;
assign addr[54873]= 931758235;
assign addr[54874]= 1000068799;
assign addr[54875]= 1067110699;
assign addr[54876]= 1132798888;
assign addr[54877]= 1197050035;
assign addr[54878]= 1259782632;
assign addr[54879]= 1320917099;
assign addr[54880]= 1380375881;
assign addr[54881]= 1438083551;
assign addr[54882]= 1493966902;
assign addr[54883]= 1547955041;
assign addr[54884]= 1599979481;
assign addr[54885]= 1649974225;
assign addr[54886]= 1697875851;
assign addr[54887]= 1743623590;
assign addr[54888]= 1787159411;
assign addr[54889]= 1828428082;
assign addr[54890]= 1867377253;
assign addr[54891]= 1903957513;
assign addr[54892]= 1938122457;
assign addr[54893]= 1969828744;
assign addr[54894]= 1999036154;
assign addr[54895]= 2025707632;
assign addr[54896]= 2049809346;
assign addr[54897]= 2071310720;
assign addr[54898]= 2090184478;
assign addr[54899]= 2106406677;
assign addr[54900]= 2119956737;
assign addr[54901]= 2130817471;
assign addr[54902]= 2138975100;
assign addr[54903]= 2144419275;
assign addr[54904]= 2147143090;
assign addr[54905]= 2147143090;
assign addr[54906]= 2144419275;
assign addr[54907]= 2138975100;
assign addr[54908]= 2130817471;
assign addr[54909]= 2119956737;
assign addr[54910]= 2106406677;
assign addr[54911]= 2090184478;
assign addr[54912]= 2071310720;
assign addr[54913]= 2049809346;
assign addr[54914]= 2025707632;
assign addr[54915]= 1999036154;
assign addr[54916]= 1969828744;
assign addr[54917]= 1938122457;
assign addr[54918]= 1903957513;
assign addr[54919]= 1867377253;
assign addr[54920]= 1828428082;
assign addr[54921]= 1787159411;
assign addr[54922]= 1743623590;
assign addr[54923]= 1697875851;
assign addr[54924]= 1649974225;
assign addr[54925]= 1599979481;
assign addr[54926]= 1547955041;
assign addr[54927]= 1493966902;
assign addr[54928]= 1438083551;
assign addr[54929]= 1380375881;
assign addr[54930]= 1320917099;
assign addr[54931]= 1259782632;
assign addr[54932]= 1197050035;
assign addr[54933]= 1132798888;
assign addr[54934]= 1067110699;
assign addr[54935]= 1000068799;
assign addr[54936]= 931758235;
assign addr[54937]= 862265664;
assign addr[54938]= 791679244;
assign addr[54939]= 720088517;
assign addr[54940]= 647584304;
assign addr[54941]= 574258580;
assign addr[54942]= 500204365;
assign addr[54943]= 425515602;
assign addr[54944]= 350287041;
assign addr[54945]= 274614114;
assign addr[54946]= 198592817;
assign addr[54947]= 122319591;
assign addr[54948]= 45891193;
assign addr[54949]= -30595422;
assign addr[54950]= -107043224;
assign addr[54951]= -183355234;
assign addr[54952]= -259434643;
assign addr[54953]= -335184940;
assign addr[54954]= -410510029;
assign addr[54955]= -485314355;
assign addr[54956]= -559503022;
assign addr[54957]= -632981917;
assign addr[54958]= -705657826;
assign addr[54959]= -777438554;
assign addr[54960]= -848233042;
assign addr[54961]= -917951481;
assign addr[54962]= -986505429;
assign addr[54963]= -1053807919;
assign addr[54964]= -1119773573;
assign addr[54965]= -1184318708;
assign addr[54966]= -1247361445;
assign addr[54967]= -1308821808;
assign addr[54968]= -1368621831;
assign addr[54969]= -1426685652;
assign addr[54970]= -1482939614;
assign addr[54971]= -1537312353;
assign addr[54972]= -1589734894;
assign addr[54973]= -1640140734;
assign addr[54974]= -1688465931;
assign addr[54975]= -1734649179;
assign addr[54976]= -1778631892;
assign addr[54977]= -1820358275;
assign addr[54978]= -1859775393;
assign addr[54979]= -1896833245;
assign addr[54980]= -1931484818;
assign addr[54981]= -1963686155;
assign addr[54982]= -1993396407;
assign addr[54983]= -2020577882;
assign addr[54984]= -2045196100;
assign addr[54985]= -2067219829;
assign addr[54986]= -2086621133;
assign addr[54987]= -2103375398;
assign addr[54988]= -2117461370;
assign addr[54989]= -2128861181;
assign addr[54990]= -2137560369;
assign addr[54991]= -2143547897;
assign addr[54992]= -2146816171;
assign addr[54993]= -2147361045;
assign addr[54994]= -2145181827;
assign addr[54995]= -2140281282;
assign addr[54996]= -2132665626;
assign addr[54997]= -2122344521;
assign addr[54998]= -2109331059;
assign addr[54999]= -2093641749;
assign addr[55000]= -2075296495;
assign addr[55001]= -2054318569;
assign addr[55002]= -2030734582;
assign addr[55003]= -2004574453;
assign addr[55004]= -1975871368;
assign addr[55005]= -1944661739;
assign addr[55006]= -1910985158;
assign addr[55007]= -1874884346;
assign addr[55008]= -1836405100;
assign addr[55009]= -1795596234;
assign addr[55010]= -1752509516;
assign addr[55011]= -1707199606;
assign addr[55012]= -1659723983;
assign addr[55013]= -1610142873;
assign addr[55014]= -1558519173;
assign addr[55015]= -1504918373;
assign addr[55016]= -1449408469;
assign addr[55017]= -1392059879;
assign addr[55018]= -1332945355;
assign addr[55019]= -1272139887;
assign addr[55020]= -1209720613;
assign addr[55021]= -1145766716;
assign addr[55022]= -1080359326;
assign addr[55023]= -1013581418;
assign addr[55024]= -945517704;
assign addr[55025]= -876254528;
assign addr[55026]= -805879757;
assign addr[55027]= -734482665;
assign addr[55028]= -662153826;
assign addr[55029]= -588984994;
assign addr[55030]= -515068990;
assign addr[55031]= -440499581;
assign addr[55032]= -365371365;
assign addr[55033]= -289779648;
assign addr[55034]= -213820322;
assign addr[55035]= -137589750;
assign addr[55036]= -61184634;
assign addr[55037]= 15298099;
assign addr[55038]= 91761426;
assign addr[55039]= 168108346;
assign addr[55040]= 244242007;
assign addr[55041]= 320065829;
assign addr[55042]= 395483624;
assign addr[55043]= 470399716;
assign addr[55044]= 544719071;
assign addr[55045]= 618347408;
assign addr[55046]= 691191324;
assign addr[55047]= 763158411;
assign addr[55048]= 834157373;
assign addr[55049]= 904098143;
assign addr[55050]= 972891995;
assign addr[55051]= 1040451659;
assign addr[55052]= 1106691431;
assign addr[55053]= 1171527280;
assign addr[55054]= 1234876957;
assign addr[55055]= 1296660098;
assign addr[55056]= 1356798326;
assign addr[55057]= 1415215352;
assign addr[55058]= 1471837070;
assign addr[55059]= 1526591649;
assign addr[55060]= 1579409630;
assign addr[55061]= 1630224009;
assign addr[55062]= 1678970324;
assign addr[55063]= 1725586737;
assign addr[55064]= 1770014111;
assign addr[55065]= 1812196087;
assign addr[55066]= 1852079154;
assign addr[55067]= 1889612716;
assign addr[55068]= 1924749160;
assign addr[55069]= 1957443913;
assign addr[55070]= 1987655498;
assign addr[55071]= 2015345591;
assign addr[55072]= 2040479063;
assign addr[55073]= 2063024031;
assign addr[55074]= 2082951896;
assign addr[55075]= 2100237377;
assign addr[55076]= 2114858546;
assign addr[55077]= 2126796855;
assign addr[55078]= 2136037160;
assign addr[55079]= 2142567738;
assign addr[55080]= 2146380306;
assign addr[55081]= 2147470025;
assign addr[55082]= 2145835515;
assign addr[55083]= 2141478848;
assign addr[55084]= 2134405552;
assign addr[55085]= 2124624598;
assign addr[55086]= 2112148396;
assign addr[55087]= 2096992772;
assign addr[55088]= 2079176953;
assign addr[55089]= 2058723538;
assign addr[55090]= 2035658475;
assign addr[55091]= 2010011024;
assign addr[55092]= 1981813720;
assign addr[55093]= 1951102334;
assign addr[55094]= 1917915825;
assign addr[55095]= 1882296293;
assign addr[55096]= 1844288924;
assign addr[55097]= 1803941934;
assign addr[55098]= 1761306505;
assign addr[55099]= 1716436725;
assign addr[55100]= 1669389513;
assign addr[55101]= 1620224553;
assign addr[55102]= 1569004214;
assign addr[55103]= 1515793473;
assign addr[55104]= 1460659832;
assign addr[55105]= 1403673233;
assign addr[55106]= 1344905966;
assign addr[55107]= 1284432584;
assign addr[55108]= 1222329801;
assign addr[55109]= 1158676398;
assign addr[55110]= 1093553126;
assign addr[55111]= 1027042599;
assign addr[55112]= 959229189;
assign addr[55113]= 890198924;
assign addr[55114]= 820039373;
assign addr[55115]= 748839539;
assign addr[55116]= 676689746;
assign addr[55117]= 603681519;
assign addr[55118]= 529907477;
assign addr[55119]= 455461206;
assign addr[55120]= 380437148;
assign addr[55121]= 304930476;
assign addr[55122]= 229036977;
assign addr[55123]= 152852926;
assign addr[55124]= 76474970;
assign addr[55125]= 0;
assign addr[55126]= -76474970;
assign addr[55127]= -152852926;
assign addr[55128]= -229036977;
assign addr[55129]= -304930476;
assign addr[55130]= -380437148;
assign addr[55131]= -455461206;
assign addr[55132]= -529907477;
assign addr[55133]= -603681519;
assign addr[55134]= -676689746;
assign addr[55135]= -748839539;
assign addr[55136]= -820039373;
assign addr[55137]= -890198924;
assign addr[55138]= -959229189;
assign addr[55139]= -1027042599;
assign addr[55140]= -1093553126;
assign addr[55141]= -1158676398;
assign addr[55142]= -1222329801;
assign addr[55143]= -1284432584;
assign addr[55144]= -1344905966;
assign addr[55145]= -1403673233;
assign addr[55146]= -1460659832;
assign addr[55147]= -1515793473;
assign addr[55148]= -1569004214;
assign addr[55149]= -1620224553;
assign addr[55150]= -1669389513;
assign addr[55151]= -1716436725;
assign addr[55152]= -1761306505;
assign addr[55153]= -1803941934;
assign addr[55154]= -1844288924;
assign addr[55155]= -1882296293;
assign addr[55156]= -1917915825;
assign addr[55157]= -1951102334;
assign addr[55158]= -1981813720;
assign addr[55159]= -2010011024;
assign addr[55160]= -2035658475;
assign addr[55161]= -2058723538;
assign addr[55162]= -2079176953;
assign addr[55163]= -2096992772;
assign addr[55164]= -2112148396;
assign addr[55165]= -2124624598;
assign addr[55166]= -2134405552;
assign addr[55167]= -2141478848;
assign addr[55168]= -2145835515;
assign addr[55169]= -2147470025;
assign addr[55170]= -2146380306;
assign addr[55171]= -2142567738;
assign addr[55172]= -2136037160;
assign addr[55173]= -2126796855;
assign addr[55174]= -2114858546;
assign addr[55175]= -2100237377;
assign addr[55176]= -2082951896;
assign addr[55177]= -2063024031;
assign addr[55178]= -2040479063;
assign addr[55179]= -2015345591;
assign addr[55180]= -1987655498;
assign addr[55181]= -1957443913;
assign addr[55182]= -1924749160;
assign addr[55183]= -1889612716;
assign addr[55184]= -1852079154;
assign addr[55185]= -1812196087;
assign addr[55186]= -1770014111;
assign addr[55187]= -1725586737;
assign addr[55188]= -1678970324;
assign addr[55189]= -1630224009;
assign addr[55190]= -1579409630;
assign addr[55191]= -1526591649;
assign addr[55192]= -1471837070;
assign addr[55193]= -1415215352;
assign addr[55194]= -1356798326;
assign addr[55195]= -1296660098;
assign addr[55196]= -1234876957;
assign addr[55197]= -1171527280;
assign addr[55198]= -1106691431;
assign addr[55199]= -1040451659;
assign addr[55200]= -972891995;
assign addr[55201]= -904098143;
assign addr[55202]= -834157373;
assign addr[55203]= -763158411;
assign addr[55204]= -691191324;
assign addr[55205]= -618347408;
assign addr[55206]= -544719071;
assign addr[55207]= -470399716;
assign addr[55208]= -395483624;
assign addr[55209]= -320065829;
assign addr[55210]= -244242007;
assign addr[55211]= -168108346;
assign addr[55212]= -91761426;
assign addr[55213]= -15298099;
assign addr[55214]= 61184634;
assign addr[55215]= 137589750;
assign addr[55216]= 213820322;
assign addr[55217]= 289779648;
assign addr[55218]= 365371365;
assign addr[55219]= 440499581;
assign addr[55220]= 515068990;
assign addr[55221]= 588984994;
assign addr[55222]= 662153826;
assign addr[55223]= 734482665;
assign addr[55224]= 805879757;
assign addr[55225]= 876254528;
assign addr[55226]= 945517704;
assign addr[55227]= 1013581418;
assign addr[55228]= 1080359326;
assign addr[55229]= 1145766716;
assign addr[55230]= 1209720613;
assign addr[55231]= 1272139887;
assign addr[55232]= 1332945355;
assign addr[55233]= 1392059879;
assign addr[55234]= 1449408469;
assign addr[55235]= 1504918373;
assign addr[55236]= 1558519173;
assign addr[55237]= 1610142873;
assign addr[55238]= 1659723983;
assign addr[55239]= 1707199606;
assign addr[55240]= 1752509516;
assign addr[55241]= 1795596234;
assign addr[55242]= 1836405100;
assign addr[55243]= 1874884346;
assign addr[55244]= 1910985158;
assign addr[55245]= 1944661739;
assign addr[55246]= 1975871368;
assign addr[55247]= 2004574453;
assign addr[55248]= 2030734582;
assign addr[55249]= 2054318569;
assign addr[55250]= 2075296495;
assign addr[55251]= 2093641749;
assign addr[55252]= 2109331059;
assign addr[55253]= 2122344521;
assign addr[55254]= 2132665626;
assign addr[55255]= 2140281282;
assign addr[55256]= 2145181827;
assign addr[55257]= 2147361045;
assign addr[55258]= 2146816171;
assign addr[55259]= 2143547897;
assign addr[55260]= 2137560369;
assign addr[55261]= 2128861181;
assign addr[55262]= 2117461370;
assign addr[55263]= 2103375398;
assign addr[55264]= 2086621133;
assign addr[55265]= 2067219829;
assign addr[55266]= 2045196100;
assign addr[55267]= 2020577882;
assign addr[55268]= 1993396407;
assign addr[55269]= 1963686155;
assign addr[55270]= 1931484818;
assign addr[55271]= 1896833245;
assign addr[55272]= 1859775393;
assign addr[55273]= 1820358275;
assign addr[55274]= 1778631892;
assign addr[55275]= 1734649179;
assign addr[55276]= 1688465931;
assign addr[55277]= 1640140734;
assign addr[55278]= 1589734894;
assign addr[55279]= 1537312353;
assign addr[55280]= 1482939614;
assign addr[55281]= 1426685652;
assign addr[55282]= 1368621831;
assign addr[55283]= 1308821808;
assign addr[55284]= 1247361445;
assign addr[55285]= 1184318708;
assign addr[55286]= 1119773573;
assign addr[55287]= 1053807919;
assign addr[55288]= 986505429;
assign addr[55289]= 917951481;
assign addr[55290]= 848233042;
assign addr[55291]= 777438554;
assign addr[55292]= 705657826;
assign addr[55293]= 632981917;
assign addr[55294]= 559503022;
assign addr[55295]= 485314355;
assign addr[55296]= 410510029;
assign addr[55297]= 335184940;
assign addr[55298]= 259434643;
assign addr[55299]= 183355234;
assign addr[55300]= 107043224;
assign addr[55301]= 30595422;
assign addr[55302]= -45891193;
assign addr[55303]= -122319591;
assign addr[55304]= -198592817;
assign addr[55305]= -274614114;
assign addr[55306]= -350287041;
assign addr[55307]= -425515602;
assign addr[55308]= -500204365;
assign addr[55309]= -574258580;
assign addr[55310]= -647584304;
assign addr[55311]= -720088517;
assign addr[55312]= -791679244;
assign addr[55313]= -862265664;
assign addr[55314]= -931758235;
assign addr[55315]= -1000068799;
assign addr[55316]= -1067110699;
assign addr[55317]= -1132798888;
assign addr[55318]= -1197050035;
assign addr[55319]= -1259782632;
assign addr[55320]= -1320917099;
assign addr[55321]= -1380375881;
assign addr[55322]= -1438083551;
assign addr[55323]= -1493966902;
assign addr[55324]= -1547955041;
assign addr[55325]= -1599979481;
assign addr[55326]= -1649974225;
assign addr[55327]= -1697875851;
assign addr[55328]= -1743623590;
assign addr[55329]= -1787159411;
assign addr[55330]= -1828428082;
assign addr[55331]= -1867377253;
assign addr[55332]= -1903957513;
assign addr[55333]= -1938122457;
assign addr[55334]= -1969828744;
assign addr[55335]= -1999036154;
assign addr[55336]= -2025707632;
assign addr[55337]= -2049809346;
assign addr[55338]= -2071310720;
assign addr[55339]= -2090184478;
assign addr[55340]= -2106406677;
assign addr[55341]= -2119956737;
assign addr[55342]= -2130817471;
assign addr[55343]= -2138975100;
assign addr[55344]= -2144419275;
assign addr[55345]= -2147143090;
assign addr[55346]= -2147143090;
assign addr[55347]= -2144419275;
assign addr[55348]= -2138975100;
assign addr[55349]= -2130817471;
assign addr[55350]= -2119956737;
assign addr[55351]= -2106406677;
assign addr[55352]= -2090184478;
assign addr[55353]= -2071310720;
assign addr[55354]= -2049809346;
assign addr[55355]= -2025707632;
assign addr[55356]= -1999036154;
assign addr[55357]= -1969828744;
assign addr[55358]= -1938122457;
assign addr[55359]= -1903957513;
assign addr[55360]= -1867377253;
assign addr[55361]= -1828428082;
assign addr[55362]= -1787159411;
assign addr[55363]= -1743623590;
assign addr[55364]= -1697875851;
assign addr[55365]= -1649974225;
assign addr[55366]= -1599979481;
assign addr[55367]= -1547955041;
assign addr[55368]= -1493966902;
assign addr[55369]= -1438083551;
assign addr[55370]= -1380375881;
assign addr[55371]= -1320917099;
assign addr[55372]= -1259782632;
assign addr[55373]= -1197050035;
assign addr[55374]= -1132798888;
assign addr[55375]= -1067110699;
assign addr[55376]= -1000068799;
assign addr[55377]= -931758235;
assign addr[55378]= -862265664;
assign addr[55379]= -791679244;
assign addr[55380]= -720088517;
assign addr[55381]= -647584304;
assign addr[55382]= -574258580;
assign addr[55383]= -500204365;
assign addr[55384]= -425515602;
assign addr[55385]= -350287041;
assign addr[55386]= -274614114;
assign addr[55387]= -198592817;
assign addr[55388]= -122319591;
assign addr[55389]= -45891193;
assign addr[55390]= 30595422;
assign addr[55391]= 107043224;
assign addr[55392]= 183355234;
assign addr[55393]= 259434643;
assign addr[55394]= 335184940;
assign addr[55395]= 410510029;
assign addr[55396]= 485314355;
assign addr[55397]= 559503022;
assign addr[55398]= 632981917;
assign addr[55399]= 705657826;
assign addr[55400]= 777438554;
assign addr[55401]= 848233042;
assign addr[55402]= 917951481;
assign addr[55403]= 986505429;
assign addr[55404]= 1053807919;
assign addr[55405]= 1119773573;
assign addr[55406]= 1184318708;
assign addr[55407]= 1247361445;
assign addr[55408]= 1308821808;
assign addr[55409]= 1368621831;
assign addr[55410]= 1426685652;
assign addr[55411]= 1482939614;
assign addr[55412]= 1537312353;
assign addr[55413]= 1589734894;
assign addr[55414]= 1640140734;
assign addr[55415]= 1688465931;
assign addr[55416]= 1734649179;
assign addr[55417]= 1778631892;
assign addr[55418]= 1820358275;
assign addr[55419]= 1859775393;
assign addr[55420]= 1896833245;
assign addr[55421]= 1931484818;
assign addr[55422]= 1963686155;
assign addr[55423]= 1993396407;
assign addr[55424]= 2020577882;
assign addr[55425]= 2045196100;
assign addr[55426]= 2067219829;
assign addr[55427]= 2086621133;
assign addr[55428]= 2103375398;
assign addr[55429]= 2117461370;
assign addr[55430]= 2128861181;
assign addr[55431]= 2137560369;
assign addr[55432]= 2143547897;
assign addr[55433]= 2146816171;
assign addr[55434]= 2147361045;
assign addr[55435]= 2145181827;
assign addr[55436]= 2140281282;
assign addr[55437]= 2132665626;
assign addr[55438]= 2122344521;
assign addr[55439]= 2109331059;
assign addr[55440]= 2093641749;
assign addr[55441]= 2075296495;
assign addr[55442]= 2054318569;
assign addr[55443]= 2030734582;
assign addr[55444]= 2004574453;
assign addr[55445]= 1975871368;
assign addr[55446]= 1944661739;
assign addr[55447]= 1910985158;
assign addr[55448]= 1874884346;
assign addr[55449]= 1836405100;
assign addr[55450]= 1795596234;
assign addr[55451]= 1752509516;
assign addr[55452]= 1707199606;
assign addr[55453]= 1659723983;
assign addr[55454]= 1610142873;
assign addr[55455]= 1558519173;
assign addr[55456]= 1504918373;
assign addr[55457]= 1449408469;
assign addr[55458]= 1392059879;
assign addr[55459]= 1332945355;
assign addr[55460]= 1272139887;
assign addr[55461]= 1209720613;
assign addr[55462]= 1145766716;
assign addr[55463]= 1080359326;
assign addr[55464]= 1013581418;
assign addr[55465]= 945517704;
assign addr[55466]= 876254528;
assign addr[55467]= 805879757;
assign addr[55468]= 734482665;
assign addr[55469]= 662153826;
assign addr[55470]= 588984994;
assign addr[55471]= 515068990;
assign addr[55472]= 440499581;
assign addr[55473]= 365371365;
assign addr[55474]= 289779648;
assign addr[55475]= 213820322;
assign addr[55476]= 137589750;
assign addr[55477]= 61184634;
assign addr[55478]= -15298099;
assign addr[55479]= -91761426;
assign addr[55480]= -168108346;
assign addr[55481]= -244242007;
assign addr[55482]= -320065829;
assign addr[55483]= -395483624;
assign addr[55484]= -470399716;
assign addr[55485]= -544719071;
assign addr[55486]= -618347408;
assign addr[55487]= -691191324;
assign addr[55488]= -763158411;
assign addr[55489]= -834157373;
assign addr[55490]= -904098143;
assign addr[55491]= -972891995;
assign addr[55492]= -1040451659;
assign addr[55493]= -1106691431;
assign addr[55494]= -1171527280;
assign addr[55495]= -1234876957;
assign addr[55496]= -1296660098;
assign addr[55497]= -1356798326;
assign addr[55498]= -1415215352;
assign addr[55499]= -1471837070;
assign addr[55500]= -1526591649;
assign addr[55501]= -1579409630;
assign addr[55502]= -1630224009;
assign addr[55503]= -1678970324;
assign addr[55504]= -1725586737;
assign addr[55505]= -1770014111;
assign addr[55506]= -1812196087;
assign addr[55507]= -1852079154;
assign addr[55508]= -1889612716;
assign addr[55509]= -1924749160;
assign addr[55510]= -1957443913;
assign addr[55511]= -1987655498;
assign addr[55512]= -2015345591;
assign addr[55513]= -2040479063;
assign addr[55514]= -2063024031;
assign addr[55515]= -2082951896;
assign addr[55516]= -2100237377;
assign addr[55517]= -2114858546;
assign addr[55518]= -2126796855;
assign addr[55519]= -2136037160;
assign addr[55520]= -2142567738;
assign addr[55521]= -2146380306;
assign addr[55522]= -2147470025;
assign addr[55523]= -2145835515;
assign addr[55524]= -2141478848;
assign addr[55525]= -2134405552;
assign addr[55526]= -2124624598;
assign addr[55527]= -2112148396;
assign addr[55528]= -2096992772;
assign addr[55529]= -2079176953;
assign addr[55530]= -2058723538;
assign addr[55531]= -2035658475;
assign addr[55532]= -2010011024;
assign addr[55533]= -1981813720;
assign addr[55534]= -1951102334;
assign addr[55535]= -1917915825;
assign addr[55536]= -1882296293;
assign addr[55537]= -1844288924;
assign addr[55538]= -1803941934;
assign addr[55539]= -1761306505;
assign addr[55540]= -1716436725;
assign addr[55541]= -1669389513;
assign addr[55542]= -1620224553;
assign addr[55543]= -1569004214;
assign addr[55544]= -1515793473;
assign addr[55545]= -1460659832;
assign addr[55546]= -1403673233;
assign addr[55547]= -1344905966;
assign addr[55548]= -1284432584;
assign addr[55549]= -1222329801;
assign addr[55550]= -1158676398;
assign addr[55551]= -1093553126;
assign addr[55552]= -1027042599;
assign addr[55553]= -959229189;
assign addr[55554]= -890198924;
assign addr[55555]= -820039373;
assign addr[55556]= -748839539;
assign addr[55557]= -676689746;
assign addr[55558]= -603681519;
assign addr[55559]= -529907477;
assign addr[55560]= -455461206;
assign addr[55561]= -380437148;
assign addr[55562]= -304930476;
assign addr[55563]= -229036977;
assign addr[55564]= -152852926;
assign addr[55565]= -76474970;
assign addr[55566]= 0;
assign addr[55567]= 76474970;
assign addr[55568]= 152852926;
assign addr[55569]= 229036977;
assign addr[55570]= 304930476;
assign addr[55571]= 380437148;
assign addr[55572]= 455461206;
assign addr[55573]= 529907477;
assign addr[55574]= 603681519;
assign addr[55575]= 676689746;
assign addr[55576]= 748839539;
assign addr[55577]= 820039373;
assign addr[55578]= 890198924;
assign addr[55579]= 959229189;
assign addr[55580]= 1027042599;
assign addr[55581]= 1093553126;
assign addr[55582]= 1158676398;
assign addr[55583]= 1222329801;
assign addr[55584]= 1284432584;
assign addr[55585]= 1344905966;
assign addr[55586]= 1403673233;
assign addr[55587]= 1460659832;
assign addr[55588]= 1515793473;
assign addr[55589]= 1569004214;
assign addr[55590]= 1620224553;
assign addr[55591]= 1669389513;
assign addr[55592]= 1716436725;
assign addr[55593]= 1761306505;
assign addr[55594]= 1803941934;
assign addr[55595]= 1844288924;
assign addr[55596]= 1882296293;
assign addr[55597]= 1917915825;
assign addr[55598]= 1951102334;
assign addr[55599]= 1981813720;
assign addr[55600]= 2010011024;
assign addr[55601]= 2035658475;
assign addr[55602]= 2058723538;
assign addr[55603]= 2079176953;
assign addr[55604]= 2096992772;
assign addr[55605]= 2112148396;
assign addr[55606]= 2124624598;
assign addr[55607]= 2134405552;
assign addr[55608]= 2141478848;
assign addr[55609]= 2145835515;
assign addr[55610]= 2147470025;
assign addr[55611]= 2146380306;
assign addr[55612]= 2142567738;
assign addr[55613]= 2136037160;
assign addr[55614]= 2126796855;
assign addr[55615]= 2114858546;
assign addr[55616]= 2100237377;
assign addr[55617]= 2082951896;
assign addr[55618]= 2063024031;
assign addr[55619]= 2040479063;
assign addr[55620]= 2015345591;
assign addr[55621]= 1987655498;
assign addr[55622]= 1957443913;
assign addr[55623]= 1924749160;
assign addr[55624]= 1889612716;
assign addr[55625]= 1852079154;
assign addr[55626]= 1812196087;
assign addr[55627]= 1770014111;
assign addr[55628]= 1725586737;
assign addr[55629]= 1678970324;
assign addr[55630]= 1630224009;
assign addr[55631]= 1579409630;
assign addr[55632]= 1526591649;
assign addr[55633]= 1471837070;
assign addr[55634]= 1415215352;
assign addr[55635]= 1356798326;
assign addr[55636]= 1296660098;
assign addr[55637]= 1234876957;
assign addr[55638]= 1171527280;
assign addr[55639]= 1106691431;
assign addr[55640]= 1040451659;
assign addr[55641]= 972891995;
assign addr[55642]= 904098143;
assign addr[55643]= 834157373;
assign addr[55644]= 763158411;
assign addr[55645]= 691191324;
assign addr[55646]= 618347408;
assign addr[55647]= 544719071;
assign addr[55648]= 470399716;
assign addr[55649]= 395483624;
assign addr[55650]= 320065829;
assign addr[55651]= 244242007;
assign addr[55652]= 168108346;
assign addr[55653]= 91761426;
assign addr[55654]= 15298099;
assign addr[55655]= -61184634;
assign addr[55656]= -137589750;
assign addr[55657]= -213820322;
assign addr[55658]= -289779648;
assign addr[55659]= -365371365;
assign addr[55660]= -440499581;
assign addr[55661]= -515068990;
assign addr[55662]= -588984994;
assign addr[55663]= -662153826;
assign addr[55664]= -734482665;
assign addr[55665]= -805879757;
assign addr[55666]= -876254528;
assign addr[55667]= -945517704;
assign addr[55668]= -1013581418;
assign addr[55669]= -1080359326;
assign addr[55670]= -1145766716;
assign addr[55671]= -1209720613;
assign addr[55672]= -1272139887;
assign addr[55673]= -1332945355;
assign addr[55674]= -1392059879;
assign addr[55675]= -1449408469;
assign addr[55676]= -1504918373;
assign addr[55677]= -1558519173;
assign addr[55678]= -1610142873;
assign addr[55679]= -1659723983;
assign addr[55680]= -1707199606;
assign addr[55681]= -1752509516;
assign addr[55682]= -1795596234;
assign addr[55683]= -1836405100;
assign addr[55684]= -1874884346;
assign addr[55685]= -1910985158;
assign addr[55686]= -1944661739;
assign addr[55687]= -1975871368;
assign addr[55688]= -2004574453;
assign addr[55689]= -2030734582;
assign addr[55690]= -2054318569;
assign addr[55691]= -2075296495;
assign addr[55692]= -2093641749;
assign addr[55693]= -2109331059;
assign addr[55694]= -2122344521;
assign addr[55695]= -2132665626;
assign addr[55696]= -2140281282;
assign addr[55697]= -2145181827;
assign addr[55698]= -2147361045;
assign addr[55699]= -2146816171;
assign addr[55700]= -2143547897;
assign addr[55701]= -2137560369;
assign addr[55702]= -2128861181;
assign addr[55703]= -2117461370;
assign addr[55704]= -2103375398;
assign addr[55705]= -2086621133;
assign addr[55706]= -2067219829;
assign addr[55707]= -2045196100;
assign addr[55708]= -2020577882;
assign addr[55709]= -1993396407;
assign addr[55710]= -1963686155;
assign addr[55711]= -1931484818;
assign addr[55712]= -1896833245;
assign addr[55713]= -1859775393;
assign addr[55714]= -1820358275;
assign addr[55715]= -1778631892;
assign addr[55716]= -1734649179;
assign addr[55717]= -1688465931;
assign addr[55718]= -1640140734;
assign addr[55719]= -1589734894;
assign addr[55720]= -1537312353;
assign addr[55721]= -1482939614;
assign addr[55722]= -1426685652;
assign addr[55723]= -1368621831;
assign addr[55724]= -1308821808;
assign addr[55725]= -1247361445;
assign addr[55726]= -1184318708;
assign addr[55727]= -1119773573;
assign addr[55728]= -1053807919;
assign addr[55729]= -986505429;
assign addr[55730]= -917951481;
assign addr[55731]= -848233042;
assign addr[55732]= -777438554;
assign addr[55733]= -705657826;
assign addr[55734]= -632981917;
assign addr[55735]= -559503022;
assign addr[55736]= -485314355;
assign addr[55737]= -410510029;
assign addr[55738]= -335184940;
assign addr[55739]= -259434643;
assign addr[55740]= -183355234;
assign addr[55741]= -107043224;
assign addr[55742]= -30595422;
assign addr[55743]= 45891193;
assign addr[55744]= 122319591;
assign addr[55745]= 198592817;
assign addr[55746]= 274614114;
assign addr[55747]= 350287041;
assign addr[55748]= 425515602;
assign addr[55749]= 500204365;
assign addr[55750]= 574258580;
assign addr[55751]= 647584304;
assign addr[55752]= 720088517;
assign addr[55753]= 791679244;
assign addr[55754]= 862265664;
assign addr[55755]= 931758235;
assign addr[55756]= 1000068799;
assign addr[55757]= 1067110699;
assign addr[55758]= 1132798888;
assign addr[55759]= 1197050035;
assign addr[55760]= 1259782632;
assign addr[55761]= 1320917099;
assign addr[55762]= 1380375881;
assign addr[55763]= 1438083551;
assign addr[55764]= 1493966902;
assign addr[55765]= 1547955041;
assign addr[55766]= 1599979481;
assign addr[55767]= 1649974225;
assign addr[55768]= 1697875851;
assign addr[55769]= 1743623590;
assign addr[55770]= 1787159411;
assign addr[55771]= 1828428082;
assign addr[55772]= 1867377253;
assign addr[55773]= 1903957513;
assign addr[55774]= 1938122457;
assign addr[55775]= 1969828744;
assign addr[55776]= 1999036154;
assign addr[55777]= 2025707632;
assign addr[55778]= 2049809346;
assign addr[55779]= 2071310720;
assign addr[55780]= 2090184478;
assign addr[55781]= 2106406677;
assign addr[55782]= 2119956737;
assign addr[55783]= 2130817471;
assign addr[55784]= 2138975100;
assign addr[55785]= 2144419275;
assign addr[55786]= 2147143090;
assign addr[55787]= 2147143090;
assign addr[55788]= 2144419275;
assign addr[55789]= 2138975100;
assign addr[55790]= 2130817471;
assign addr[55791]= 2119956737;
assign addr[55792]= 2106406677;
assign addr[55793]= 2090184478;
assign addr[55794]= 2071310720;
assign addr[55795]= 2049809346;
assign addr[55796]= 2025707632;
assign addr[55797]= 1999036154;
assign addr[55798]= 1969828744;
assign addr[55799]= 1938122457;
assign addr[55800]= 1903957513;
assign addr[55801]= 1867377253;
assign addr[55802]= 1828428082;
assign addr[55803]= 1787159411;
assign addr[55804]= 1743623590;
assign addr[55805]= 1697875851;
assign addr[55806]= 1649974225;
assign addr[55807]= 1599979481;
assign addr[55808]= 1547955041;
assign addr[55809]= 1493966902;
assign addr[55810]= 1438083551;
assign addr[55811]= 1380375881;
assign addr[55812]= 1320917099;
assign addr[55813]= 1259782632;
assign addr[55814]= 1197050035;
assign addr[55815]= 1132798888;
assign addr[55816]= 1067110699;
assign addr[55817]= 1000068799;
assign addr[55818]= 931758235;
assign addr[55819]= 862265664;
assign addr[55820]= 791679244;
assign addr[55821]= 720088517;
assign addr[55822]= 647584304;
assign addr[55823]= 574258580;
assign addr[55824]= 500204365;
assign addr[55825]= 425515602;
assign addr[55826]= 350287041;
assign addr[55827]= 274614114;
assign addr[55828]= 198592817;
assign addr[55829]= 122319591;
assign addr[55830]= 45891193;
assign addr[55831]= -30595422;
assign addr[55832]= -107043224;
assign addr[55833]= -183355234;
assign addr[55834]= -259434643;
assign addr[55835]= -335184940;
assign addr[55836]= -410510029;
assign addr[55837]= -485314355;
assign addr[55838]= -559503022;
assign addr[55839]= -632981917;
assign addr[55840]= -705657826;
assign addr[55841]= -777438554;
assign addr[55842]= -848233042;
assign addr[55843]= -917951481;
assign addr[55844]= -986505429;
assign addr[55845]= -1053807919;
assign addr[55846]= -1119773573;
assign addr[55847]= -1184318708;
assign addr[55848]= -1247361445;
assign addr[55849]= -1308821808;
assign addr[55850]= -1368621831;
assign addr[55851]= -1426685652;
assign addr[55852]= -1482939614;
assign addr[55853]= -1537312353;
assign addr[55854]= -1589734894;
assign addr[55855]= -1640140734;
assign addr[55856]= -1688465931;
assign addr[55857]= -1734649179;
assign addr[55858]= -1778631892;
assign addr[55859]= -1820358275;
assign addr[55860]= -1859775393;
assign addr[55861]= -1896833245;
assign addr[55862]= -1931484818;
assign addr[55863]= -1963686155;
assign addr[55864]= -1993396407;
assign addr[55865]= -2020577882;
assign addr[55866]= -2045196100;
assign addr[55867]= -2067219829;
assign addr[55868]= -2086621133;
assign addr[55869]= -2103375398;
assign addr[55870]= -2117461370;
assign addr[55871]= -2128861181;
assign addr[55872]= -2137560369;
assign addr[55873]= -2143547897;
assign addr[55874]= -2146816171;
assign addr[55875]= -2147361045;
assign addr[55876]= -2145181827;
assign addr[55877]= -2140281282;
assign addr[55878]= -2132665626;
assign addr[55879]= -2122344521;
assign addr[55880]= -2109331059;
assign addr[55881]= -2093641749;
assign addr[55882]= -2075296495;
assign addr[55883]= -2054318569;
assign addr[55884]= -2030734582;
assign addr[55885]= -2004574453;
assign addr[55886]= -1975871368;
assign addr[55887]= -1944661739;
assign addr[55888]= -1910985158;
assign addr[55889]= -1874884346;
assign addr[55890]= -1836405100;
assign addr[55891]= -1795596234;
assign addr[55892]= -1752509516;
assign addr[55893]= -1707199606;
assign addr[55894]= -1659723983;
assign addr[55895]= -1610142873;
assign addr[55896]= -1558519173;
assign addr[55897]= -1504918373;
assign addr[55898]= -1449408469;
assign addr[55899]= -1392059879;
assign addr[55900]= -1332945355;
assign addr[55901]= -1272139887;
assign addr[55902]= -1209720613;
assign addr[55903]= -1145766716;
assign addr[55904]= -1080359326;
assign addr[55905]= -1013581418;
assign addr[55906]= -945517704;
assign addr[55907]= -876254528;
assign addr[55908]= -805879757;
assign addr[55909]= -734482665;
assign addr[55910]= -662153826;
assign addr[55911]= -588984994;
assign addr[55912]= -515068990;
assign addr[55913]= -440499581;
assign addr[55914]= -365371365;
assign addr[55915]= -289779648;
assign addr[55916]= -213820322;
assign addr[55917]= -137589750;
assign addr[55918]= -61184634;
assign addr[55919]= 15298099;
assign addr[55920]= 91761426;
assign addr[55921]= 168108346;
assign addr[55922]= 244242007;
assign addr[55923]= 320065829;
assign addr[55924]= 395483624;
assign addr[55925]= 470399716;
assign addr[55926]= 544719071;
assign addr[55927]= 618347408;
assign addr[55928]= 691191324;
assign addr[55929]= 763158411;
assign addr[55930]= 834157373;
assign addr[55931]= 904098143;
assign addr[55932]= 972891995;
assign addr[55933]= 1040451659;
assign addr[55934]= 1106691431;
assign addr[55935]= 1171527280;
assign addr[55936]= 1234876957;
assign addr[55937]= 1296660098;
assign addr[55938]= 1356798326;
assign addr[55939]= 1415215352;
assign addr[55940]= 1471837070;
assign addr[55941]= 1526591649;
assign addr[55942]= 1579409630;
assign addr[55943]= 1630224009;
assign addr[55944]= 1678970324;
assign addr[55945]= 1725586737;
assign addr[55946]= 1770014111;
assign addr[55947]= 1812196087;
assign addr[55948]= 1852079154;
assign addr[55949]= 1889612716;
assign addr[55950]= 1924749160;
assign addr[55951]= 1957443913;
assign addr[55952]= 1987655498;
assign addr[55953]= 2015345591;
assign addr[55954]= 2040479063;
assign addr[55955]= 2063024031;
assign addr[55956]= 2082951896;
assign addr[55957]= 2100237377;
assign addr[55958]= 2114858546;
assign addr[55959]= 2126796855;
assign addr[55960]= 2136037160;
assign addr[55961]= 2142567738;
assign addr[55962]= 2146380306;
assign addr[55963]= 2147470025;
assign addr[55964]= 2145835515;
assign addr[55965]= 2141478848;
assign addr[55966]= 2134405552;
assign addr[55967]= 2124624598;
assign addr[55968]= 2112148396;
assign addr[55969]= 2096992772;
assign addr[55970]= 2079176953;
assign addr[55971]= 2058723538;
assign addr[55972]= 2035658475;
assign addr[55973]= 2010011024;
assign addr[55974]= 1981813720;
assign addr[55975]= 1951102334;
assign addr[55976]= 1917915825;
assign addr[55977]= 1882296293;
assign addr[55978]= 1844288924;
assign addr[55979]= 1803941934;
assign addr[55980]= 1761306505;
assign addr[55981]= 1716436725;
assign addr[55982]= 1669389513;
assign addr[55983]= 1620224553;
assign addr[55984]= 1569004214;
assign addr[55985]= 1515793473;
assign addr[55986]= 1460659832;
assign addr[55987]= 1403673233;
assign addr[55988]= 1344905966;
assign addr[55989]= 1284432584;
assign addr[55990]= 1222329801;
assign addr[55991]= 1158676398;
assign addr[55992]= 1093553126;
assign addr[55993]= 1027042599;
assign addr[55994]= 959229189;
assign addr[55995]= 890198924;
assign addr[55996]= 820039373;
assign addr[55997]= 748839539;
assign addr[55998]= 676689746;
assign addr[55999]= 603681519;
assign addr[56000]= 529907477;
assign addr[56001]= 455461206;
assign addr[56002]= 380437148;
assign addr[56003]= 304930476;
assign addr[56004]= 229036977;
assign addr[56005]= 152852926;
assign addr[56006]= 76474970;
assign addr[56007]= 0;
assign addr[56008]= -76474970;
assign addr[56009]= -152852926;
assign addr[56010]= -229036977;
assign addr[56011]= -304930476;
assign addr[56012]= -380437148;
assign addr[56013]= -455461206;
assign addr[56014]= -529907477;
assign addr[56015]= -603681519;
assign addr[56016]= -676689746;
assign addr[56017]= -748839539;
assign addr[56018]= -820039373;
assign addr[56019]= -890198924;
assign addr[56020]= -959229189;
assign addr[56021]= -1027042599;
assign addr[56022]= -1093553126;
assign addr[56023]= -1158676398;
assign addr[56024]= -1222329801;
assign addr[56025]= -1284432584;
assign addr[56026]= -1344905966;
assign addr[56027]= -1403673233;
assign addr[56028]= -1460659832;
assign addr[56029]= -1515793473;
assign addr[56030]= -1569004214;
assign addr[56031]= -1620224553;
assign addr[56032]= -1669389513;
assign addr[56033]= -1716436725;
assign addr[56034]= -1761306505;
assign addr[56035]= -1803941934;
assign addr[56036]= -1844288924;
assign addr[56037]= -1882296293;
assign addr[56038]= -1917915825;
assign addr[56039]= -1951102334;
assign addr[56040]= -1981813720;
assign addr[56041]= -2010011024;
assign addr[56042]= -2035658475;
assign addr[56043]= -2058723538;
assign addr[56044]= -2079176953;
assign addr[56045]= -2096992772;
assign addr[56046]= -2112148396;
assign addr[56047]= -2124624598;
assign addr[56048]= -2134405552;
assign addr[56049]= -2141478848;
assign addr[56050]= -2145835515;
assign addr[56051]= -2147470025;
assign addr[56052]= -2146380306;
assign addr[56053]= -2142567738;
assign addr[56054]= -2136037160;
assign addr[56055]= -2126796855;
assign addr[56056]= -2114858546;
assign addr[56057]= -2100237377;
assign addr[56058]= -2082951896;
assign addr[56059]= -2063024031;
assign addr[56060]= -2040479063;
assign addr[56061]= -2015345591;
assign addr[56062]= -1987655498;
assign addr[56063]= -1957443913;
assign addr[56064]= -1924749160;
assign addr[56065]= -1889612716;
assign addr[56066]= -1852079154;
assign addr[56067]= -1812196087;
assign addr[56068]= -1770014111;
assign addr[56069]= -1725586737;
assign addr[56070]= -1678970324;
assign addr[56071]= -1630224009;
assign addr[56072]= -1579409630;
assign addr[56073]= -1526591649;
assign addr[56074]= -1471837070;
assign addr[56075]= -1415215352;
assign addr[56076]= -1356798326;
assign addr[56077]= -1296660098;
assign addr[56078]= -1234876957;
assign addr[56079]= -1171527280;
assign addr[56080]= -1106691431;
assign addr[56081]= -1040451659;
assign addr[56082]= -972891995;
assign addr[56083]= -904098143;
assign addr[56084]= -834157373;
assign addr[56085]= -763158411;
assign addr[56086]= -691191324;
assign addr[56087]= -618347408;
assign addr[56088]= -544719071;
assign addr[56089]= -470399716;
assign addr[56090]= -395483624;
assign addr[56091]= -320065829;
assign addr[56092]= -244242007;
assign addr[56093]= -168108346;
assign addr[56094]= -91761426;
assign addr[56095]= -15298099;
assign addr[56096]= 61184634;
assign addr[56097]= 137589750;
assign addr[56098]= 213820322;
assign addr[56099]= 289779648;
assign addr[56100]= 365371365;
assign addr[56101]= 440499581;
assign addr[56102]= 515068990;
assign addr[56103]= 588984994;
assign addr[56104]= 662153826;
assign addr[56105]= 734482665;
assign addr[56106]= 805879757;
assign addr[56107]= 876254528;
assign addr[56108]= 945517704;
assign addr[56109]= 1013581418;
assign addr[56110]= 1080359326;
assign addr[56111]= 1145766716;
assign addr[56112]= 1209720613;
assign addr[56113]= 1272139887;
assign addr[56114]= 1332945355;
assign addr[56115]= 1392059879;
assign addr[56116]= 1449408469;
assign addr[56117]= 1504918373;
assign addr[56118]= 1558519173;
assign addr[56119]= 1610142873;
assign addr[56120]= 1659723983;
assign addr[56121]= 1707199606;
assign addr[56122]= 1752509516;
assign addr[56123]= 1795596234;
assign addr[56124]= 1836405100;
assign addr[56125]= 1874884346;
assign addr[56126]= 1910985158;
assign addr[56127]= 1944661739;
assign addr[56128]= 1975871368;
assign addr[56129]= 2004574453;
assign addr[56130]= 2030734582;
assign addr[56131]= 2054318569;
assign addr[56132]= 2075296495;
assign addr[56133]= 2093641749;
assign addr[56134]= 2109331059;
assign addr[56135]= 2122344521;
assign addr[56136]= 2132665626;
assign addr[56137]= 2140281282;
assign addr[56138]= 2145181827;
assign addr[56139]= 2147361045;
assign addr[56140]= 2146816171;
assign addr[56141]= 2143547897;
assign addr[56142]= 2137560369;
assign addr[56143]= 2128861181;
assign addr[56144]= 2117461370;
assign addr[56145]= 2103375398;
assign addr[56146]= 2086621133;
assign addr[56147]= 2067219829;
assign addr[56148]= 2045196100;
assign addr[56149]= 2020577882;
assign addr[56150]= 1993396407;
assign addr[56151]= 1963686155;
assign addr[56152]= 1931484818;
assign addr[56153]= 1896833245;
assign addr[56154]= 1859775393;
assign addr[56155]= 1820358275;
assign addr[56156]= 1778631892;
assign addr[56157]= 1734649179;
assign addr[56158]= 1688465931;
assign addr[56159]= 1640140734;
assign addr[56160]= 1589734894;
assign addr[56161]= 1537312353;
assign addr[56162]= 1482939614;
assign addr[56163]= 1426685652;
assign addr[56164]= 1368621831;
assign addr[56165]= 1308821808;
assign addr[56166]= 1247361445;
assign addr[56167]= 1184318708;
assign addr[56168]= 1119773573;
assign addr[56169]= 1053807919;
assign addr[56170]= 986505429;
assign addr[56171]= 917951481;
assign addr[56172]= 848233042;
assign addr[56173]= 777438554;
assign addr[56174]= 705657826;
assign addr[56175]= 632981917;
assign addr[56176]= 559503022;
assign addr[56177]= 485314355;
assign addr[56178]= 410510029;
assign addr[56179]= 335184940;
assign addr[56180]= 259434643;
assign addr[56181]= 183355234;
assign addr[56182]= 107043224;
assign addr[56183]= 30595422;
assign addr[56184]= -45891193;
assign addr[56185]= -122319591;
assign addr[56186]= -198592817;
assign addr[56187]= -274614114;
assign addr[56188]= -350287041;
assign addr[56189]= -425515602;
assign addr[56190]= -500204365;
assign addr[56191]= -574258580;
assign addr[56192]= -647584304;
assign addr[56193]= -720088517;
assign addr[56194]= -791679244;
assign addr[56195]= -862265664;
assign addr[56196]= -931758235;
assign addr[56197]= -1000068799;
assign addr[56198]= -1067110699;
assign addr[56199]= -1132798888;
assign addr[56200]= -1197050035;
assign addr[56201]= -1259782632;
assign addr[56202]= -1320917099;
assign addr[56203]= -1380375881;
assign addr[56204]= -1438083551;
assign addr[56205]= -1493966902;
assign addr[56206]= -1547955041;
assign addr[56207]= -1599979481;
assign addr[56208]= -1649974225;
assign addr[56209]= -1697875851;
assign addr[56210]= -1743623590;
assign addr[56211]= -1787159411;
assign addr[56212]= -1828428082;
assign addr[56213]= -1867377253;
assign addr[56214]= -1903957513;
assign addr[56215]= -1938122457;
assign addr[56216]= -1969828744;
assign addr[56217]= -1999036154;
assign addr[56218]= -2025707632;
assign addr[56219]= -2049809346;
assign addr[56220]= -2071310720;
assign addr[56221]= -2090184478;
assign addr[56222]= -2106406677;
assign addr[56223]= -2119956737;
assign addr[56224]= -2130817471;
assign addr[56225]= -2138975100;
assign addr[56226]= -2144419275;
assign addr[56227]= -2147143090;
assign addr[56228]= -2147143090;
assign addr[56229]= -2144419275;
assign addr[56230]= -2138975100;
assign addr[56231]= -2130817471;
assign addr[56232]= -2119956737;
assign addr[56233]= -2106406677;
assign addr[56234]= -2090184478;
assign addr[56235]= -2071310720;
assign addr[56236]= -2049809346;
assign addr[56237]= -2025707632;
assign addr[56238]= -1999036154;
assign addr[56239]= -1969828744;
assign addr[56240]= -1938122457;
assign addr[56241]= -1903957513;
assign addr[56242]= -1867377253;
assign addr[56243]= -1828428082;
assign addr[56244]= -1787159411;
assign addr[56245]= -1743623590;
assign addr[56246]= -1697875851;
assign addr[56247]= -1649974225;
assign addr[56248]= -1599979481;
assign addr[56249]= -1547955041;
assign addr[56250]= -1493966902;
assign addr[56251]= -1438083551;
assign addr[56252]= -1380375881;
assign addr[56253]= -1320917099;
assign addr[56254]= -1259782632;
assign addr[56255]= -1197050035;
assign addr[56256]= -1132798888;
assign addr[56257]= -1067110699;
assign addr[56258]= -1000068799;
assign addr[56259]= -931758235;
assign addr[56260]= -862265664;
assign addr[56261]= -791679244;
assign addr[56262]= -720088517;
assign addr[56263]= -647584304;
assign addr[56264]= -574258580;
assign addr[56265]= -500204365;
assign addr[56266]= -425515602;
assign addr[56267]= -350287041;
assign addr[56268]= -274614114;
assign addr[56269]= -198592817;
assign addr[56270]= -122319591;
assign addr[56271]= -45891193;
assign addr[56272]= 30595422;
assign addr[56273]= 107043224;
assign addr[56274]= 183355234;
assign addr[56275]= 259434643;
assign addr[56276]= 335184940;
assign addr[56277]= 410510029;
assign addr[56278]= 485314355;
assign addr[56279]= 559503022;
assign addr[56280]= 632981917;
assign addr[56281]= 705657826;
assign addr[56282]= 777438554;
assign addr[56283]= 848233042;
assign addr[56284]= 917951481;
assign addr[56285]= 986505429;
assign addr[56286]= 1053807919;
assign addr[56287]= 1119773573;
assign addr[56288]= 1184318708;
assign addr[56289]= 1247361445;
assign addr[56290]= 1308821808;
assign addr[56291]= 1368621831;
assign addr[56292]= 1426685652;
assign addr[56293]= 1482939614;
assign addr[56294]= 1537312353;
assign addr[56295]= 1589734894;
assign addr[56296]= 1640140734;
assign addr[56297]= 1688465931;
assign addr[56298]= 1734649179;
assign addr[56299]= 1778631892;
assign addr[56300]= 1820358275;
assign addr[56301]= 1859775393;
assign addr[56302]= 1896833245;
assign addr[56303]= 1931484818;
assign addr[56304]= 1963686155;
assign addr[56305]= 1993396407;
assign addr[56306]= 2020577882;
assign addr[56307]= 2045196100;
assign addr[56308]= 2067219829;
assign addr[56309]= 2086621133;
assign addr[56310]= 2103375398;
assign addr[56311]= 2117461370;
assign addr[56312]= 2128861181;
assign addr[56313]= 2137560369;
assign addr[56314]= 2143547897;
assign addr[56315]= 2146816171;
assign addr[56316]= 2147361045;
assign addr[56317]= 2145181827;
assign addr[56318]= 2140281282;
assign addr[56319]= 2132665626;
assign addr[56320]= 2122344521;
assign addr[56321]= 2109331059;
assign addr[56322]= 2093641749;
assign addr[56323]= 2075296495;
assign addr[56324]= 2054318569;
assign addr[56325]= 2030734582;
assign addr[56326]= 2004574453;
assign addr[56327]= 1975871368;
assign addr[56328]= 1944661739;
assign addr[56329]= 1910985158;
assign addr[56330]= 1874884346;
assign addr[56331]= 1836405100;
assign addr[56332]= 1795596234;
assign addr[56333]= 1752509516;
assign addr[56334]= 1707199606;
assign addr[56335]= 1659723983;
assign addr[56336]= 1610142873;
assign addr[56337]= 1558519173;
assign addr[56338]= 1504918373;
assign addr[56339]= 1449408469;
assign addr[56340]= 1392059879;
assign addr[56341]= 1332945355;
assign addr[56342]= 1272139887;
assign addr[56343]= 1209720613;
assign addr[56344]= 1145766716;
assign addr[56345]= 1080359326;
assign addr[56346]= 1013581418;
assign addr[56347]= 945517704;
assign addr[56348]= 876254528;
assign addr[56349]= 805879757;
assign addr[56350]= 734482665;
assign addr[56351]= 662153826;
assign addr[56352]= 588984994;
assign addr[56353]= 515068990;
assign addr[56354]= 440499581;
assign addr[56355]= 365371365;
assign addr[56356]= 289779648;
assign addr[56357]= 213820322;
assign addr[56358]= 137589750;
assign addr[56359]= 61184634;
assign addr[56360]= -15298099;
assign addr[56361]= -91761426;
assign addr[56362]= -168108346;
assign addr[56363]= -244242007;
assign addr[56364]= -320065829;
assign addr[56365]= -395483624;
assign addr[56366]= -470399716;
assign addr[56367]= -544719071;
assign addr[56368]= -618347408;
assign addr[56369]= -691191324;
assign addr[56370]= -763158411;
assign addr[56371]= -834157373;
assign addr[56372]= -904098143;
assign addr[56373]= -972891995;
assign addr[56374]= -1040451659;
assign addr[56375]= -1106691431;
assign addr[56376]= -1171527280;
assign addr[56377]= -1234876957;
assign addr[56378]= -1296660098;
assign addr[56379]= -1356798326;
assign addr[56380]= -1415215352;
assign addr[56381]= -1471837070;
assign addr[56382]= -1526591649;
assign addr[56383]= -1579409630;
assign addr[56384]= -1630224009;
assign addr[56385]= -1678970324;
assign addr[56386]= -1725586737;
assign addr[56387]= -1770014111;
assign addr[56388]= -1812196087;
assign addr[56389]= -1852079154;
assign addr[56390]= -1889612716;
assign addr[56391]= -1924749160;
assign addr[56392]= -1957443913;
assign addr[56393]= -1987655498;
assign addr[56394]= -2015345591;
assign addr[56395]= -2040479063;
assign addr[56396]= -2063024031;
assign addr[56397]= -2082951896;
assign addr[56398]= -2100237377;
assign addr[56399]= -2114858546;
assign addr[56400]= -2126796855;
assign addr[56401]= -2136037160;
assign addr[56402]= -2142567738;
assign addr[56403]= -2146380306;
assign addr[56404]= -2147470025;
assign addr[56405]= -2145835515;
assign addr[56406]= -2141478848;
assign addr[56407]= -2134405552;
assign addr[56408]= -2124624598;
assign addr[56409]= -2112148396;
assign addr[56410]= -2096992772;
assign addr[56411]= -2079176953;
assign addr[56412]= -2058723538;
assign addr[56413]= -2035658475;
assign addr[56414]= -2010011024;
assign addr[56415]= -1981813720;
assign addr[56416]= -1951102334;
assign addr[56417]= -1917915825;
assign addr[56418]= -1882296293;
assign addr[56419]= -1844288924;
assign addr[56420]= -1803941934;
assign addr[56421]= -1761306505;
assign addr[56422]= -1716436725;
assign addr[56423]= -1669389513;
assign addr[56424]= -1620224553;
assign addr[56425]= -1569004214;
assign addr[56426]= -1515793473;
assign addr[56427]= -1460659832;
assign addr[56428]= -1403673233;
assign addr[56429]= -1344905966;
assign addr[56430]= -1284432584;
assign addr[56431]= -1222329801;
assign addr[56432]= -1158676398;
assign addr[56433]= -1093553126;
assign addr[56434]= -1027042599;
assign addr[56435]= -959229189;
assign addr[56436]= -890198924;
assign addr[56437]= -820039373;
assign addr[56438]= -748839539;
assign addr[56439]= -676689746;
assign addr[56440]= -603681519;
assign addr[56441]= -529907477;
assign addr[56442]= -455461206;
assign addr[56443]= -380437148;
assign addr[56444]= -304930476;
assign addr[56445]= -229036977;
assign addr[56446]= -152852926;
assign addr[56447]= -76474970;
assign addr[56448]= 0;
assign addr[56449]= 76474970;
assign addr[56450]= 152852926;
assign addr[56451]= 229036977;
assign addr[56452]= 304930476;
assign addr[56453]= 380437148;
assign addr[56454]= 455461206;
assign addr[56455]= 529907477;
assign addr[56456]= 603681519;
assign addr[56457]= 676689746;
assign addr[56458]= 748839539;
assign addr[56459]= 820039373;
assign addr[56460]= 890198924;
assign addr[56461]= 959229189;
assign addr[56462]= 1027042599;
assign addr[56463]= 1093553126;
assign addr[56464]= 1158676398;
assign addr[56465]= 1222329801;
assign addr[56466]= 1284432584;
assign addr[56467]= 1344905966;
assign addr[56468]= 1403673233;
assign addr[56469]= 1460659832;
assign addr[56470]= 1515793473;
assign addr[56471]= 1569004214;
assign addr[56472]= 1620224553;
assign addr[56473]= 1669389513;
assign addr[56474]= 1716436725;
assign addr[56475]= 1761306505;
assign addr[56476]= 1803941934;
assign addr[56477]= 1844288924;
assign addr[56478]= 1882296293;
assign addr[56479]= 1917915825;
assign addr[56480]= 1951102334;
assign addr[56481]= 1981813720;
assign addr[56482]= 2010011024;
assign addr[56483]= 2035658475;
assign addr[56484]= 2058723538;
assign addr[56485]= 2079176953;
assign addr[56486]= 2096992772;
assign addr[56487]= 2112148396;
assign addr[56488]= 2124624598;
assign addr[56489]= 2134405552;
assign addr[56490]= 2141478848;
assign addr[56491]= 2145835515;
assign addr[56492]= 2147470025;
assign addr[56493]= 2146380306;
assign addr[56494]= 2142567738;
assign addr[56495]= 2136037160;
assign addr[56496]= 2126796855;
assign addr[56497]= 2114858546;
assign addr[56498]= 2100237377;
assign addr[56499]= 2082951896;
assign addr[56500]= 2063024031;
assign addr[56501]= 2040479063;
assign addr[56502]= 2015345591;
assign addr[56503]= 1987655498;
assign addr[56504]= 1957443913;
assign addr[56505]= 1924749160;
assign addr[56506]= 1889612716;
assign addr[56507]= 1852079154;
assign addr[56508]= 1812196087;
assign addr[56509]= 1770014111;
assign addr[56510]= 1725586737;
assign addr[56511]= 1678970324;
assign addr[56512]= 1630224009;
assign addr[56513]= 1579409630;
assign addr[56514]= 1526591649;
assign addr[56515]= 1471837070;
assign addr[56516]= 1415215352;
assign addr[56517]= 1356798326;
assign addr[56518]= 1296660098;
assign addr[56519]= 1234876957;
assign addr[56520]= 1171527280;
assign addr[56521]= 1106691431;
assign addr[56522]= 1040451659;
assign addr[56523]= 972891995;
assign addr[56524]= 904098143;
assign addr[56525]= 834157373;
assign addr[56526]= 763158411;
assign addr[56527]= 691191324;
assign addr[56528]= 618347408;
assign addr[56529]= 544719071;
assign addr[56530]= 470399716;
assign addr[56531]= 395483624;
assign addr[56532]= 320065829;
assign addr[56533]= 244242007;
assign addr[56534]= 168108346;
assign addr[56535]= 91761426;
assign addr[56536]= 15298099;
assign addr[56537]= -61184634;
assign addr[56538]= -137589750;
assign addr[56539]= -213820322;
assign addr[56540]= -289779648;
assign addr[56541]= -365371365;
assign addr[56542]= -440499581;
assign addr[56543]= -515068990;
assign addr[56544]= -588984994;
assign addr[56545]= -662153826;
assign addr[56546]= -734482665;
assign addr[56547]= -805879757;
assign addr[56548]= -876254528;
assign addr[56549]= -945517704;
assign addr[56550]= -1013581418;
assign addr[56551]= -1080359326;
assign addr[56552]= -1145766716;
assign addr[56553]= -1209720613;
assign addr[56554]= -1272139887;
assign addr[56555]= -1332945355;
assign addr[56556]= -1392059879;
assign addr[56557]= -1449408469;
assign addr[56558]= -1504918373;
assign addr[56559]= -1558519173;
assign addr[56560]= -1610142873;
assign addr[56561]= -1659723983;
assign addr[56562]= -1707199606;
assign addr[56563]= -1752509516;
assign addr[56564]= -1795596234;
assign addr[56565]= -1836405100;
assign addr[56566]= -1874884346;
assign addr[56567]= -1910985158;
assign addr[56568]= -1944661739;
assign addr[56569]= -1975871368;
assign addr[56570]= -2004574453;
assign addr[56571]= -2030734582;
assign addr[56572]= -2054318569;
assign addr[56573]= -2075296495;
assign addr[56574]= -2093641749;
assign addr[56575]= -2109331059;
assign addr[56576]= -2122344521;
assign addr[56577]= -2132665626;
assign addr[56578]= -2140281282;
assign addr[56579]= -2145181827;
assign addr[56580]= -2147361045;
assign addr[56581]= -2146816171;
assign addr[56582]= -2143547897;
assign addr[56583]= -2137560369;
assign addr[56584]= -2128861181;
assign addr[56585]= -2117461370;
assign addr[56586]= -2103375398;
assign addr[56587]= -2086621133;
assign addr[56588]= -2067219829;
assign addr[56589]= -2045196100;
assign addr[56590]= -2020577882;
assign addr[56591]= -1993396407;
assign addr[56592]= -1963686155;
assign addr[56593]= -1931484818;
assign addr[56594]= -1896833245;
assign addr[56595]= -1859775393;
assign addr[56596]= -1820358275;
assign addr[56597]= -1778631892;
assign addr[56598]= -1734649179;
assign addr[56599]= -1688465931;
assign addr[56600]= -1640140734;
assign addr[56601]= -1589734894;
assign addr[56602]= -1537312353;
assign addr[56603]= -1482939614;
assign addr[56604]= -1426685652;
assign addr[56605]= -1368621831;
assign addr[56606]= -1308821808;
assign addr[56607]= -1247361445;
assign addr[56608]= -1184318708;
assign addr[56609]= -1119773573;
assign addr[56610]= -1053807919;
assign addr[56611]= -986505429;
assign addr[56612]= -917951481;
assign addr[56613]= -848233042;
assign addr[56614]= -777438554;
assign addr[56615]= -705657826;
assign addr[56616]= -632981917;
assign addr[56617]= -559503022;
assign addr[56618]= -485314355;
assign addr[56619]= -410510029;
assign addr[56620]= -335184940;
assign addr[56621]= -259434643;
assign addr[56622]= -183355234;
assign addr[56623]= -107043224;
assign addr[56624]= -30595422;
assign addr[56625]= 45891193;
assign addr[56626]= 122319591;
assign addr[56627]= 198592817;
assign addr[56628]= 274614114;
assign addr[56629]= 350287041;
assign addr[56630]= 425515602;
assign addr[56631]= 500204365;
assign addr[56632]= 574258580;
assign addr[56633]= 647584304;
assign addr[56634]= 720088517;
assign addr[56635]= 791679244;
assign addr[56636]= 862265664;
assign addr[56637]= 931758235;
assign addr[56638]= 1000068799;
assign addr[56639]= 1067110699;
assign addr[56640]= 1132798888;
assign addr[56641]= 1197050035;
assign addr[56642]= 1259782632;
assign addr[56643]= 1320917099;
assign addr[56644]= 1380375881;
assign addr[56645]= 1438083551;
assign addr[56646]= 1493966902;
assign addr[56647]= 1547955041;
assign addr[56648]= 1599979481;
assign addr[56649]= 1649974225;
assign addr[56650]= 1697875851;
assign addr[56651]= 1743623590;
assign addr[56652]= 1787159411;
assign addr[56653]= 1828428082;
assign addr[56654]= 1867377253;
assign addr[56655]= 1903957513;
assign addr[56656]= 1938122457;
assign addr[56657]= 1969828744;
assign addr[56658]= 1999036154;
assign addr[56659]= 2025707632;
assign addr[56660]= 2049809346;
assign addr[56661]= 2071310720;
assign addr[56662]= 2090184478;
assign addr[56663]= 2106406677;
assign addr[56664]= 2119956737;
assign addr[56665]= 2130817471;
assign addr[56666]= 2138975100;
assign addr[56667]= 2144419275;
assign addr[56668]= 2147143090;
assign addr[56669]= 2147143090;
assign addr[56670]= 2144419275;
assign addr[56671]= 2138975100;
assign addr[56672]= 2130817471;
assign addr[56673]= 2119956737;
assign addr[56674]= 2106406677;
assign addr[56675]= 2090184478;
assign addr[56676]= 2071310720;
assign addr[56677]= 2049809346;
assign addr[56678]= 2025707632;
assign addr[56679]= 1999036154;
assign addr[56680]= 1969828744;
assign addr[56681]= 1938122457;
assign addr[56682]= 1903957513;
assign addr[56683]= 1867377253;
assign addr[56684]= 1828428082;
assign addr[56685]= 1787159411;
assign addr[56686]= 1743623590;
assign addr[56687]= 1697875851;
assign addr[56688]= 1649974225;
assign addr[56689]= 1599979481;
assign addr[56690]= 1547955041;
assign addr[56691]= 1493966902;
assign addr[56692]= 1438083551;
assign addr[56693]= 1380375881;
assign addr[56694]= 1320917099;
assign addr[56695]= 1259782632;
assign addr[56696]= 1197050035;
assign addr[56697]= 1132798888;
assign addr[56698]= 1067110699;
assign addr[56699]= 1000068799;
assign addr[56700]= 931758235;
assign addr[56701]= 862265664;
assign addr[56702]= 791679244;
assign addr[56703]= 720088517;
assign addr[56704]= 647584304;
assign addr[56705]= 574258580;
assign addr[56706]= 500204365;
assign addr[56707]= 425515602;
assign addr[56708]= 350287041;
assign addr[56709]= 274614114;
assign addr[56710]= 198592817;
assign addr[56711]= 122319591;
assign addr[56712]= 45891193;
assign addr[56713]= -30595422;
assign addr[56714]= -107043224;
assign addr[56715]= -183355234;
assign addr[56716]= -259434643;
assign addr[56717]= -335184940;
assign addr[56718]= -410510029;
assign addr[56719]= -485314355;
assign addr[56720]= -559503022;
assign addr[56721]= -632981917;
assign addr[56722]= -705657826;
assign addr[56723]= -777438554;
assign addr[56724]= -848233042;
assign addr[56725]= -917951481;
assign addr[56726]= -986505429;
assign addr[56727]= -1053807919;
assign addr[56728]= -1119773573;
assign addr[56729]= -1184318708;
assign addr[56730]= -1247361445;
assign addr[56731]= -1308821808;
assign addr[56732]= -1368621831;
assign addr[56733]= -1426685652;
assign addr[56734]= -1482939614;
assign addr[56735]= -1537312353;
assign addr[56736]= -1589734894;
assign addr[56737]= -1640140734;
assign addr[56738]= -1688465931;
assign addr[56739]= -1734649179;
assign addr[56740]= -1778631892;
assign addr[56741]= -1820358275;
assign addr[56742]= -1859775393;
assign addr[56743]= -1896833245;
assign addr[56744]= -1931484818;
assign addr[56745]= -1963686155;
assign addr[56746]= -1993396407;
assign addr[56747]= -2020577882;
assign addr[56748]= -2045196100;
assign addr[56749]= -2067219829;
assign addr[56750]= -2086621133;
assign addr[56751]= -2103375398;
assign addr[56752]= -2117461370;
assign addr[56753]= -2128861181;
assign addr[56754]= -2137560369;
assign addr[56755]= -2143547897;
assign addr[56756]= -2146816171;
assign addr[56757]= -2147361045;
assign addr[56758]= -2145181827;
assign addr[56759]= -2140281282;
assign addr[56760]= -2132665626;
assign addr[56761]= -2122344521;
assign addr[56762]= -2109331059;
assign addr[56763]= -2093641749;
assign addr[56764]= -2075296495;
assign addr[56765]= -2054318569;
assign addr[56766]= -2030734582;
assign addr[56767]= -2004574453;
assign addr[56768]= -1975871368;
assign addr[56769]= -1944661739;
assign addr[56770]= -1910985158;
assign addr[56771]= -1874884346;
assign addr[56772]= -1836405100;
assign addr[56773]= -1795596234;
assign addr[56774]= -1752509516;
assign addr[56775]= -1707199606;
assign addr[56776]= -1659723983;
assign addr[56777]= -1610142873;
assign addr[56778]= -1558519173;
assign addr[56779]= -1504918373;
assign addr[56780]= -1449408469;
assign addr[56781]= -1392059879;
assign addr[56782]= -1332945355;
assign addr[56783]= -1272139887;
assign addr[56784]= -1209720613;
assign addr[56785]= -1145766716;
assign addr[56786]= -1080359326;
assign addr[56787]= -1013581418;
assign addr[56788]= -945517704;
assign addr[56789]= -876254528;
assign addr[56790]= -805879757;
assign addr[56791]= -734482665;
assign addr[56792]= -662153826;
assign addr[56793]= -588984994;
assign addr[56794]= -515068990;
assign addr[56795]= -440499581;
assign addr[56796]= -365371365;
assign addr[56797]= -289779648;
assign addr[56798]= -213820322;
assign addr[56799]= -137589750;
assign addr[56800]= -61184634;
assign addr[56801]= 15298099;
assign addr[56802]= 91761426;
assign addr[56803]= 168108346;
assign addr[56804]= 244242007;
assign addr[56805]= 320065829;
assign addr[56806]= 395483624;
assign addr[56807]= 470399716;
assign addr[56808]= 544719071;
assign addr[56809]= 618347408;
assign addr[56810]= 691191324;
assign addr[56811]= 763158411;
assign addr[56812]= 834157373;
assign addr[56813]= 904098143;
assign addr[56814]= 972891995;
assign addr[56815]= 1040451659;
assign addr[56816]= 1106691431;
assign addr[56817]= 1171527280;
assign addr[56818]= 1234876957;
assign addr[56819]= 1296660098;
assign addr[56820]= 1356798326;
assign addr[56821]= 1415215352;
assign addr[56822]= 1471837070;
assign addr[56823]= 1526591649;
assign addr[56824]= 1579409630;
assign addr[56825]= 1630224009;
assign addr[56826]= 1678970324;
assign addr[56827]= 1725586737;
assign addr[56828]= 1770014111;
assign addr[56829]= 1812196087;
assign addr[56830]= 1852079154;
assign addr[56831]= 1889612716;
assign addr[56832]= 1924749160;
assign addr[56833]= 1957443913;
assign addr[56834]= 1987655498;
assign addr[56835]= 2015345591;
assign addr[56836]= 2040479063;
assign addr[56837]= 2063024031;
assign addr[56838]= 2082951896;
assign addr[56839]= 2100237377;
assign addr[56840]= 2114858546;
assign addr[56841]= 2126796855;
assign addr[56842]= 2136037160;
assign addr[56843]= 2142567738;
assign addr[56844]= 2146380306;
assign addr[56845]= 2147470025;
assign addr[56846]= 2145835515;
assign addr[56847]= 2141478848;
assign addr[56848]= 2134405552;
assign addr[56849]= 2124624598;
assign addr[56850]= 2112148396;
assign addr[56851]= 2096992772;
assign addr[56852]= 2079176953;
assign addr[56853]= 2058723538;
assign addr[56854]= 2035658475;
assign addr[56855]= 2010011024;
assign addr[56856]= 1981813720;
assign addr[56857]= 1951102334;
assign addr[56858]= 1917915825;
assign addr[56859]= 1882296293;
assign addr[56860]= 1844288924;
assign addr[56861]= 1803941934;
assign addr[56862]= 1761306505;
assign addr[56863]= 1716436725;
assign addr[56864]= 1669389513;
assign addr[56865]= 1620224553;
assign addr[56866]= 1569004214;
assign addr[56867]= 1515793473;
assign addr[56868]= 1460659832;
assign addr[56869]= 1403673233;
assign addr[56870]= 1344905966;
assign addr[56871]= 1284432584;
assign addr[56872]= 1222329801;
assign addr[56873]= 1158676398;
assign addr[56874]= 1093553126;
assign addr[56875]= 1027042599;
assign addr[56876]= 959229189;
assign addr[56877]= 890198924;
assign addr[56878]= 820039373;
assign addr[56879]= 748839539;
assign addr[56880]= 676689746;
assign addr[56881]= 603681519;
assign addr[56882]= 529907477;
assign addr[56883]= 455461206;
assign addr[56884]= 380437148;
assign addr[56885]= 304930476;
assign addr[56886]= 229036977;
assign addr[56887]= 152852926;
assign addr[56888]= 76474970;
assign addr[56889]= 0;
assign addr[56890]= -76474970;
assign addr[56891]= -152852926;
assign addr[56892]= -229036977;
assign addr[56893]= -304930476;
assign addr[56894]= -380437148;
assign addr[56895]= -455461206;
assign addr[56896]= -529907477;
assign addr[56897]= -603681519;
assign addr[56898]= -676689746;
assign addr[56899]= -748839539;
assign addr[56900]= -820039373;
assign addr[56901]= -890198924;
assign addr[56902]= -959229189;
assign addr[56903]= -1027042599;
assign addr[56904]= -1093553126;
assign addr[56905]= -1158676398;
assign addr[56906]= -1222329801;
assign addr[56907]= -1284432584;
assign addr[56908]= -1344905966;
assign addr[56909]= -1403673233;
assign addr[56910]= -1460659832;
assign addr[56911]= -1515793473;
assign addr[56912]= -1569004214;
assign addr[56913]= -1620224553;
assign addr[56914]= -1669389513;
assign addr[56915]= -1716436725;
assign addr[56916]= -1761306505;
assign addr[56917]= -1803941934;
assign addr[56918]= -1844288924;
assign addr[56919]= -1882296293;
assign addr[56920]= -1917915825;
assign addr[56921]= -1951102334;
assign addr[56922]= -1981813720;
assign addr[56923]= -2010011024;
assign addr[56924]= -2035658475;
assign addr[56925]= -2058723538;
assign addr[56926]= -2079176953;
assign addr[56927]= -2096992772;
assign addr[56928]= -2112148396;
assign addr[56929]= -2124624598;
assign addr[56930]= -2134405552;
assign addr[56931]= -2141478848;
assign addr[56932]= -2145835515;
assign addr[56933]= -2147470025;
assign addr[56934]= -2146380306;
assign addr[56935]= -2142567738;
assign addr[56936]= -2136037160;
assign addr[56937]= -2126796855;
assign addr[56938]= -2114858546;
assign addr[56939]= -2100237377;
assign addr[56940]= -2082951896;
assign addr[56941]= -2063024031;
assign addr[56942]= -2040479063;
assign addr[56943]= -2015345591;
assign addr[56944]= -1987655498;
assign addr[56945]= -1957443913;
assign addr[56946]= -1924749160;
assign addr[56947]= -1889612716;
assign addr[56948]= -1852079154;
assign addr[56949]= -1812196087;
assign addr[56950]= -1770014111;
assign addr[56951]= -1725586737;
assign addr[56952]= -1678970324;
assign addr[56953]= -1630224009;
assign addr[56954]= -1579409630;
assign addr[56955]= -1526591649;
assign addr[56956]= -1471837070;
assign addr[56957]= -1415215352;
assign addr[56958]= -1356798326;
assign addr[56959]= -1296660098;
assign addr[56960]= -1234876957;
assign addr[56961]= -1171527280;
assign addr[56962]= -1106691431;
assign addr[56963]= -1040451659;
assign addr[56964]= -972891995;
assign addr[56965]= -904098143;
assign addr[56966]= -834157373;
assign addr[56967]= -763158411;
assign addr[56968]= -691191324;
assign addr[56969]= -618347408;
assign addr[56970]= -544719071;
assign addr[56971]= -470399716;
assign addr[56972]= -395483624;
assign addr[56973]= -320065829;
assign addr[56974]= -244242007;
assign addr[56975]= -168108346;
assign addr[56976]= -91761426;
assign addr[56977]= -15298099;
assign addr[56978]= 61184634;
assign addr[56979]= 137589750;
assign addr[56980]= 213820322;
assign addr[56981]= 289779648;
assign addr[56982]= 365371365;
assign addr[56983]= 440499581;
assign addr[56984]= 515068990;
assign addr[56985]= 588984994;
assign addr[56986]= 662153826;
assign addr[56987]= 734482665;
assign addr[56988]= 805879757;
assign addr[56989]= 876254528;
assign addr[56990]= 945517704;
assign addr[56991]= 1013581418;
assign addr[56992]= 1080359326;
assign addr[56993]= 1145766716;
assign addr[56994]= 1209720613;
assign addr[56995]= 1272139887;
assign addr[56996]= 1332945355;
assign addr[56997]= 1392059879;
assign addr[56998]= 1449408469;
assign addr[56999]= 1504918373;
assign addr[57000]= 1558519173;
assign addr[57001]= 1610142873;
assign addr[57002]= 1659723983;
assign addr[57003]= 1707199606;
assign addr[57004]= 1752509516;
assign addr[57005]= 1795596234;
assign addr[57006]= 1836405100;
assign addr[57007]= 1874884346;
assign addr[57008]= 1910985158;
assign addr[57009]= 1944661739;
assign addr[57010]= 1975871368;
assign addr[57011]= 2004574453;
assign addr[57012]= 2030734582;
assign addr[57013]= 2054318569;
assign addr[57014]= 2075296495;
assign addr[57015]= 2093641749;
assign addr[57016]= 2109331059;
assign addr[57017]= 2122344521;
assign addr[57018]= 2132665626;
assign addr[57019]= 2140281282;
assign addr[57020]= 2145181827;
assign addr[57021]= 2147361045;
assign addr[57022]= 2146816171;
assign addr[57023]= 2143547897;
assign addr[57024]= 2137560369;
assign addr[57025]= 2128861181;
assign addr[57026]= 2117461370;
assign addr[57027]= 2103375398;
assign addr[57028]= 2086621133;
assign addr[57029]= 2067219829;
assign addr[57030]= 2045196100;
assign addr[57031]= 2020577882;
assign addr[57032]= 1993396407;
assign addr[57033]= 1963686155;
assign addr[57034]= 1931484818;
assign addr[57035]= 1896833245;
assign addr[57036]= 1859775393;
assign addr[57037]= 1820358275;
assign addr[57038]= 1778631892;
assign addr[57039]= 1734649179;
assign addr[57040]= 1688465931;
assign addr[57041]= 1640140734;
assign addr[57042]= 1589734894;
assign addr[57043]= 1537312353;
assign addr[57044]= 1482939614;
assign addr[57045]= 1426685652;
assign addr[57046]= 1368621831;
assign addr[57047]= 1308821808;
assign addr[57048]= 1247361445;
assign addr[57049]= 1184318708;
assign addr[57050]= 1119773573;
assign addr[57051]= 1053807919;
assign addr[57052]= 986505429;
assign addr[57053]= 917951481;
assign addr[57054]= 848233042;
assign addr[57055]= 777438554;
assign addr[57056]= 705657826;
assign addr[57057]= 632981917;
assign addr[57058]= 559503022;
assign addr[57059]= 485314355;
assign addr[57060]= 410510029;
assign addr[57061]= 335184940;
assign addr[57062]= 259434643;
assign addr[57063]= 183355234;
assign addr[57064]= 107043224;
assign addr[57065]= 30595422;
assign addr[57066]= -45891193;
assign addr[57067]= -122319591;
assign addr[57068]= -198592817;
assign addr[57069]= -274614114;
assign addr[57070]= -350287041;
assign addr[57071]= -425515602;
assign addr[57072]= -500204365;
assign addr[57073]= -574258580;
assign addr[57074]= -647584304;
assign addr[57075]= -720088517;
assign addr[57076]= -791679244;
assign addr[57077]= -862265664;
assign addr[57078]= -931758235;
assign addr[57079]= -1000068799;
assign addr[57080]= -1067110699;
assign addr[57081]= -1132798888;
assign addr[57082]= -1197050035;
assign addr[57083]= -1259782632;
assign addr[57084]= -1320917099;
assign addr[57085]= -1380375881;
assign addr[57086]= -1438083551;
assign addr[57087]= -1493966902;
assign addr[57088]= -1547955041;
assign addr[57089]= -1599979481;
assign addr[57090]= -1649974225;
assign addr[57091]= -1697875851;
assign addr[57092]= -1743623590;
assign addr[57093]= -1787159411;
assign addr[57094]= -1828428082;
assign addr[57095]= -1867377253;
assign addr[57096]= -1903957513;
assign addr[57097]= -1938122457;
assign addr[57098]= -1969828744;
assign addr[57099]= -1999036154;
assign addr[57100]= -2025707632;
assign addr[57101]= -2049809346;
assign addr[57102]= -2071310720;
assign addr[57103]= -2090184478;
assign addr[57104]= -2106406677;
assign addr[57105]= -2119956737;
assign addr[57106]= -2130817471;
assign addr[57107]= -2138975100;
assign addr[57108]= -2144419275;
assign addr[57109]= -2147143090;
assign addr[57110]= -2147143090;
assign addr[57111]= -2144419275;
assign addr[57112]= -2138975100;
assign addr[57113]= -2130817471;
assign addr[57114]= -2119956737;
assign addr[57115]= -2106406677;
assign addr[57116]= -2090184478;
assign addr[57117]= -2071310720;
assign addr[57118]= -2049809346;
assign addr[57119]= -2025707632;
assign addr[57120]= -1999036154;
assign addr[57121]= -1969828744;
assign addr[57122]= -1938122457;
assign addr[57123]= -1903957513;
assign addr[57124]= -1867377253;
assign addr[57125]= -1828428082;
assign addr[57126]= -1787159411;
assign addr[57127]= -1743623590;
assign addr[57128]= -1697875851;
assign addr[57129]= -1649974225;
assign addr[57130]= -1599979481;
assign addr[57131]= -1547955041;
assign addr[57132]= -1493966902;
assign addr[57133]= -1438083551;
assign addr[57134]= -1380375881;
assign addr[57135]= -1320917099;
assign addr[57136]= -1259782632;
assign addr[57137]= -1197050035;
assign addr[57138]= -1132798888;
assign addr[57139]= -1067110699;
assign addr[57140]= -1000068799;
assign addr[57141]= -931758235;
assign addr[57142]= -862265664;
assign addr[57143]= -791679244;
assign addr[57144]= -720088517;
assign addr[57145]= -647584304;
assign addr[57146]= -574258580;
assign addr[57147]= -500204365;
assign addr[57148]= -425515602;
assign addr[57149]= -350287041;
assign addr[57150]= -274614114;
assign addr[57151]= -198592817;
assign addr[57152]= -122319591;
assign addr[57153]= -45891193;
assign addr[57154]= 30595422;
assign addr[57155]= 107043224;
assign addr[57156]= 183355234;
assign addr[57157]= 259434643;
assign addr[57158]= 335184940;
assign addr[57159]= 410510029;
assign addr[57160]= 485314355;
assign addr[57161]= 559503022;
assign addr[57162]= 632981917;
assign addr[57163]= 705657826;
assign addr[57164]= 777438554;
assign addr[57165]= 848233042;
assign addr[57166]= 917951481;
assign addr[57167]= 986505429;
assign addr[57168]= 1053807919;
assign addr[57169]= 1119773573;
assign addr[57170]= 1184318708;
assign addr[57171]= 1247361445;
assign addr[57172]= 1308821808;
assign addr[57173]= 1368621831;
assign addr[57174]= 1426685652;
assign addr[57175]= 1482939614;
assign addr[57176]= 1537312353;
assign addr[57177]= 1589734894;
assign addr[57178]= 1640140734;
assign addr[57179]= 1688465931;
assign addr[57180]= 1734649179;
assign addr[57181]= 1778631892;
assign addr[57182]= 1820358275;
assign addr[57183]= 1859775393;
assign addr[57184]= 1896833245;
assign addr[57185]= 1931484818;
assign addr[57186]= 1963686155;
assign addr[57187]= 1993396407;
assign addr[57188]= 2020577882;
assign addr[57189]= 2045196100;
assign addr[57190]= 2067219829;
assign addr[57191]= 2086621133;
assign addr[57192]= 2103375398;
assign addr[57193]= 2117461370;
assign addr[57194]= 2128861181;
assign addr[57195]= 2137560369;
assign addr[57196]= 2143547897;
assign addr[57197]= 2146816171;
assign addr[57198]= 2147361045;
assign addr[57199]= 2145181827;
assign addr[57200]= 2140281282;
assign addr[57201]= 2132665626;
assign addr[57202]= 2122344521;
assign addr[57203]= 2109331059;
assign addr[57204]= 2093641749;
assign addr[57205]= 2075296495;
assign addr[57206]= 2054318569;
assign addr[57207]= 2030734582;
assign addr[57208]= 2004574453;
assign addr[57209]= 1975871368;
assign addr[57210]= 1944661739;
assign addr[57211]= 1910985158;
assign addr[57212]= 1874884346;
assign addr[57213]= 1836405100;
assign addr[57214]= 1795596234;
assign addr[57215]= 1752509516;
assign addr[57216]= 1707199606;
assign addr[57217]= 1659723983;
assign addr[57218]= 1610142873;
assign addr[57219]= 1558519173;
assign addr[57220]= 1504918373;
assign addr[57221]= 1449408469;
assign addr[57222]= 1392059879;
assign addr[57223]= 1332945355;
assign addr[57224]= 1272139887;
assign addr[57225]= 1209720613;
assign addr[57226]= 1145766716;
assign addr[57227]= 1080359326;
assign addr[57228]= 1013581418;
assign addr[57229]= 945517704;
assign addr[57230]= 876254528;
assign addr[57231]= 805879757;
assign addr[57232]= 734482665;
assign addr[57233]= 662153826;
assign addr[57234]= 588984994;
assign addr[57235]= 515068990;
assign addr[57236]= 440499581;
assign addr[57237]= 365371365;
assign addr[57238]= 289779648;
assign addr[57239]= 213820322;
assign addr[57240]= 137589750;
assign addr[57241]= 61184634;
assign addr[57242]= -15298099;
assign addr[57243]= -91761426;
assign addr[57244]= -168108346;
assign addr[57245]= -244242007;
assign addr[57246]= -320065829;
assign addr[57247]= -395483624;
assign addr[57248]= -470399716;
assign addr[57249]= -544719071;
assign addr[57250]= -618347408;
assign addr[57251]= -691191324;
assign addr[57252]= -763158411;
assign addr[57253]= -834157373;
assign addr[57254]= -904098143;
assign addr[57255]= -972891995;
assign addr[57256]= -1040451659;
assign addr[57257]= -1106691431;
assign addr[57258]= -1171527280;
assign addr[57259]= -1234876957;
assign addr[57260]= -1296660098;
assign addr[57261]= -1356798326;
assign addr[57262]= -1415215352;
assign addr[57263]= -1471837070;
assign addr[57264]= -1526591649;
assign addr[57265]= -1579409630;
assign addr[57266]= -1630224009;
assign addr[57267]= -1678970324;
assign addr[57268]= -1725586737;
assign addr[57269]= -1770014111;
assign addr[57270]= -1812196087;
assign addr[57271]= -1852079154;
assign addr[57272]= -1889612716;
assign addr[57273]= -1924749160;
assign addr[57274]= -1957443913;
assign addr[57275]= -1987655498;
assign addr[57276]= -2015345591;
assign addr[57277]= -2040479063;
assign addr[57278]= -2063024031;
assign addr[57279]= -2082951896;
assign addr[57280]= -2100237377;
assign addr[57281]= -2114858546;
assign addr[57282]= -2126796855;
assign addr[57283]= -2136037160;
assign addr[57284]= -2142567738;
assign addr[57285]= -2146380306;
assign addr[57286]= -2147470025;
assign addr[57287]= -2145835515;
assign addr[57288]= -2141478848;
assign addr[57289]= -2134405552;
assign addr[57290]= -2124624598;
assign addr[57291]= -2112148396;
assign addr[57292]= -2096992772;
assign addr[57293]= -2079176953;
assign addr[57294]= -2058723538;
assign addr[57295]= -2035658475;
assign addr[57296]= -2010011024;
assign addr[57297]= -1981813720;
assign addr[57298]= -1951102334;
assign addr[57299]= -1917915825;
assign addr[57300]= -1882296293;
assign addr[57301]= -1844288924;
assign addr[57302]= -1803941934;
assign addr[57303]= -1761306505;
assign addr[57304]= -1716436725;
assign addr[57305]= -1669389513;
assign addr[57306]= -1620224553;
assign addr[57307]= -1569004214;
assign addr[57308]= -1515793473;
assign addr[57309]= -1460659832;
assign addr[57310]= -1403673233;
assign addr[57311]= -1344905966;
assign addr[57312]= -1284432584;
assign addr[57313]= -1222329801;
assign addr[57314]= -1158676398;
assign addr[57315]= -1093553126;
assign addr[57316]= -1027042599;
assign addr[57317]= -959229189;
assign addr[57318]= -890198924;
assign addr[57319]= -820039373;
assign addr[57320]= -748839539;
assign addr[57321]= -676689746;
assign addr[57322]= -603681519;
assign addr[57323]= -529907477;
assign addr[57324]= -455461206;
assign addr[57325]= -380437148;
assign addr[57326]= -304930476;
assign addr[57327]= -229036977;
assign addr[57328]= -152852926;
assign addr[57329]= -76474970;
assign addr[57330]= 0;
assign addr[57331]= 76474970;
assign addr[57332]= 152852926;
assign addr[57333]= 229036977;
assign addr[57334]= 304930476;
assign addr[57335]= 380437148;
assign addr[57336]= 455461206;
assign addr[57337]= 529907477;
assign addr[57338]= 603681519;
assign addr[57339]= 676689746;
assign addr[57340]= 748839539;
assign addr[57341]= 820039373;
assign addr[57342]= 890198924;
assign addr[57343]= 959229189;
assign addr[57344]= 1027042599;
assign addr[57345]= 1093553126;
assign addr[57346]= 1158676398;
assign addr[57347]= 1222329801;
assign addr[57348]= 1284432584;
assign addr[57349]= 1344905966;
assign addr[57350]= 1403673233;
assign addr[57351]= 1460659832;
assign addr[57352]= 1515793473;
assign addr[57353]= 1569004214;
assign addr[57354]= 1620224553;
assign addr[57355]= 1669389513;
assign addr[57356]= 1716436725;
assign addr[57357]= 1761306505;
assign addr[57358]= 1803941934;
assign addr[57359]= 1844288924;
assign addr[57360]= 1882296293;
assign addr[57361]= 1917915825;
assign addr[57362]= 1951102334;
assign addr[57363]= 1981813720;
assign addr[57364]= 2010011024;
assign addr[57365]= 2035658475;
assign addr[57366]= 2058723538;
assign addr[57367]= 2079176953;
assign addr[57368]= 2096992772;
assign addr[57369]= 2112148396;
assign addr[57370]= 2124624598;
assign addr[57371]= 2134405552;
assign addr[57372]= 2141478848;
assign addr[57373]= 2145835515;
assign addr[57374]= 2147470025;
assign addr[57375]= 2146380306;
assign addr[57376]= 2142567738;
assign addr[57377]= 2136037160;
assign addr[57378]= 2126796855;
assign addr[57379]= 2114858546;
assign addr[57380]= 2100237377;
assign addr[57381]= 2082951896;
assign addr[57382]= 2063024031;
assign addr[57383]= 2040479063;
assign addr[57384]= 2015345591;
assign addr[57385]= 1987655498;
assign addr[57386]= 1957443913;
assign addr[57387]= 1924749160;
assign addr[57388]= 1889612716;
assign addr[57389]= 1852079154;
assign addr[57390]= 1812196087;
assign addr[57391]= 1770014111;
assign addr[57392]= 1725586737;
assign addr[57393]= 1678970324;
assign addr[57394]= 1630224009;
assign addr[57395]= 1579409630;
assign addr[57396]= 1526591649;
assign addr[57397]= 1471837070;
assign addr[57398]= 1415215352;
assign addr[57399]= 1356798326;
assign addr[57400]= 1296660098;
assign addr[57401]= 1234876957;
assign addr[57402]= 1171527280;
assign addr[57403]= 1106691431;
assign addr[57404]= 1040451659;
assign addr[57405]= 972891995;
assign addr[57406]= 904098143;
assign addr[57407]= 834157373;
assign addr[57408]= 763158411;
assign addr[57409]= 691191324;
assign addr[57410]= 618347408;
assign addr[57411]= 544719071;
assign addr[57412]= 470399716;
assign addr[57413]= 395483624;
assign addr[57414]= 320065829;
assign addr[57415]= 244242007;
assign addr[57416]= 168108346;
assign addr[57417]= 91761426;
assign addr[57418]= 15298099;
assign addr[57419]= -61184634;
assign addr[57420]= -137589750;
assign addr[57421]= -213820322;
assign addr[57422]= -289779648;
assign addr[57423]= -365371365;
assign addr[57424]= -440499581;
assign addr[57425]= -515068990;
assign addr[57426]= -588984994;
assign addr[57427]= -662153826;
assign addr[57428]= -734482665;
assign addr[57429]= -805879757;
assign addr[57430]= -876254528;
assign addr[57431]= -945517704;
assign addr[57432]= -1013581418;
assign addr[57433]= -1080359326;
assign addr[57434]= -1145766716;
assign addr[57435]= -1209720613;
assign addr[57436]= -1272139887;
assign addr[57437]= -1332945355;
assign addr[57438]= -1392059879;
assign addr[57439]= -1449408469;
assign addr[57440]= -1504918373;
assign addr[57441]= -1558519173;
assign addr[57442]= -1610142873;
assign addr[57443]= -1659723983;
assign addr[57444]= -1707199606;
assign addr[57445]= -1752509516;
assign addr[57446]= -1795596234;
assign addr[57447]= -1836405100;
assign addr[57448]= -1874884346;
assign addr[57449]= -1910985158;
assign addr[57450]= -1944661739;
assign addr[57451]= -1975871368;
assign addr[57452]= -2004574453;
assign addr[57453]= -2030734582;
assign addr[57454]= -2054318569;
assign addr[57455]= -2075296495;
assign addr[57456]= -2093641749;
assign addr[57457]= -2109331059;
assign addr[57458]= -2122344521;
assign addr[57459]= -2132665626;
assign addr[57460]= -2140281282;
assign addr[57461]= -2145181827;
assign addr[57462]= -2147361045;
assign addr[57463]= -2146816171;
assign addr[57464]= -2143547897;
assign addr[57465]= -2137560369;
assign addr[57466]= -2128861181;
assign addr[57467]= -2117461370;
assign addr[57468]= -2103375398;
assign addr[57469]= -2086621133;
assign addr[57470]= -2067219829;
assign addr[57471]= -2045196100;
assign addr[57472]= -2020577882;
assign addr[57473]= -1993396407;
assign addr[57474]= -1963686155;
assign addr[57475]= -1931484818;
assign addr[57476]= -1896833245;
assign addr[57477]= -1859775393;
assign addr[57478]= -1820358275;
assign addr[57479]= -1778631892;
assign addr[57480]= -1734649179;
assign addr[57481]= -1688465931;
assign addr[57482]= -1640140734;
assign addr[57483]= -1589734894;
assign addr[57484]= -1537312353;
assign addr[57485]= -1482939614;
assign addr[57486]= -1426685652;
assign addr[57487]= -1368621831;
assign addr[57488]= -1308821808;
assign addr[57489]= -1247361445;
assign addr[57490]= -1184318708;
assign addr[57491]= -1119773573;
assign addr[57492]= -1053807919;
assign addr[57493]= -986505429;
assign addr[57494]= -917951481;
assign addr[57495]= -848233042;
assign addr[57496]= -777438554;
assign addr[57497]= -705657826;
assign addr[57498]= -632981917;
assign addr[57499]= -559503022;
assign addr[57500]= -485314355;
assign addr[57501]= -410510029;
assign addr[57502]= -335184940;
assign addr[57503]= -259434643;
assign addr[57504]= -183355234;
assign addr[57505]= -107043224;
assign addr[57506]= -30595422;
assign addr[57507]= 45891193;
assign addr[57508]= 122319591;
assign addr[57509]= 198592817;
assign addr[57510]= 274614114;
assign addr[57511]= 350287041;
assign addr[57512]= 425515602;
assign addr[57513]= 500204365;
assign addr[57514]= 574258580;
assign addr[57515]= 647584304;
assign addr[57516]= 720088517;
assign addr[57517]= 791679244;
assign addr[57518]= 862265664;
assign addr[57519]= 931758235;
assign addr[57520]= 1000068799;
assign addr[57521]= 1067110699;
assign addr[57522]= 1132798888;
assign addr[57523]= 1197050035;
assign addr[57524]= 1259782632;
assign addr[57525]= 1320917099;
assign addr[57526]= 1380375881;
assign addr[57527]= 1438083551;
assign addr[57528]= 1493966902;
assign addr[57529]= 1547955041;
assign addr[57530]= 1599979481;
assign addr[57531]= 1649974225;
assign addr[57532]= 1697875851;
assign addr[57533]= 1743623590;
assign addr[57534]= 1787159411;
assign addr[57535]= 1828428082;
assign addr[57536]= 1867377253;
assign addr[57537]= 1903957513;
assign addr[57538]= 1938122457;
assign addr[57539]= 1969828744;
assign addr[57540]= 1999036154;
assign addr[57541]= 2025707632;
assign addr[57542]= 2049809346;
assign addr[57543]= 2071310720;
assign addr[57544]= 2090184478;
assign addr[57545]= 2106406677;
assign addr[57546]= 2119956737;
assign addr[57547]= 2130817471;
assign addr[57548]= 2138975100;
assign addr[57549]= 2144419275;
assign addr[57550]= 2147143090;
assign addr[57551]= 2147143090;
assign addr[57552]= 2144419275;
assign addr[57553]= 2138975100;
assign addr[57554]= 2130817471;
assign addr[57555]= 2119956737;
assign addr[57556]= 2106406677;
assign addr[57557]= 2090184478;
assign addr[57558]= 2071310720;
assign addr[57559]= 2049809346;
assign addr[57560]= 2025707632;
assign addr[57561]= 1999036154;
assign addr[57562]= 1969828744;
assign addr[57563]= 1938122457;
assign addr[57564]= 1903957513;
assign addr[57565]= 1867377253;
assign addr[57566]= 1828428082;
assign addr[57567]= 1787159411;
assign addr[57568]= 1743623590;
assign addr[57569]= 1697875851;
assign addr[57570]= 1649974225;
assign addr[57571]= 1599979481;
assign addr[57572]= 1547955041;
assign addr[57573]= 1493966902;
assign addr[57574]= 1438083551;
assign addr[57575]= 1380375881;
assign addr[57576]= 1320917099;
assign addr[57577]= 1259782632;
assign addr[57578]= 1197050035;
assign addr[57579]= 1132798888;
assign addr[57580]= 1067110699;
assign addr[57581]= 1000068799;
assign addr[57582]= 931758235;
assign addr[57583]= 862265664;
assign addr[57584]= 791679244;
assign addr[57585]= 720088517;
assign addr[57586]= 647584304;
assign addr[57587]= 574258580;
assign addr[57588]= 500204365;
assign addr[57589]= 425515602;
assign addr[57590]= 350287041;
assign addr[57591]= 274614114;
assign addr[57592]= 198592817;
assign addr[57593]= 122319591;
assign addr[57594]= 45891193;
assign addr[57595]= -30595422;
assign addr[57596]= -107043224;
assign addr[57597]= -183355234;
assign addr[57598]= -259434643;
assign addr[57599]= -335184940;
assign addr[57600]= -410510029;
assign addr[57601]= -485314355;
assign addr[57602]= -559503022;
assign addr[57603]= -632981917;
assign addr[57604]= -705657826;
assign addr[57605]= -777438554;
assign addr[57606]= -848233042;
assign addr[57607]= -917951481;
assign addr[57608]= -986505429;
assign addr[57609]= -1053807919;
assign addr[57610]= -1119773573;
assign addr[57611]= -1184318708;
assign addr[57612]= -1247361445;
assign addr[57613]= -1308821808;
assign addr[57614]= -1368621831;
assign addr[57615]= -1426685652;
assign addr[57616]= -1482939614;
assign addr[57617]= -1537312353;
assign addr[57618]= -1589734894;
assign addr[57619]= -1640140734;
assign addr[57620]= -1688465931;
assign addr[57621]= -1734649179;
assign addr[57622]= -1778631892;
assign addr[57623]= -1820358275;
assign addr[57624]= -1859775393;
assign addr[57625]= -1896833245;
assign addr[57626]= -1931484818;
assign addr[57627]= -1963686155;
assign addr[57628]= -1993396407;
assign addr[57629]= -2020577882;
assign addr[57630]= -2045196100;
assign addr[57631]= -2067219829;
assign addr[57632]= -2086621133;
assign addr[57633]= -2103375398;
assign addr[57634]= -2117461370;
assign addr[57635]= -2128861181;
assign addr[57636]= -2137560369;
assign addr[57637]= -2143547897;
assign addr[57638]= -2146816171;
assign addr[57639]= -2147361045;
assign addr[57640]= -2145181827;
assign addr[57641]= -2140281282;
assign addr[57642]= -2132665626;
assign addr[57643]= -2122344521;
assign addr[57644]= -2109331059;
assign addr[57645]= -2093641749;
assign addr[57646]= -2075296495;
assign addr[57647]= -2054318569;
assign addr[57648]= -2030734582;
assign addr[57649]= -2004574453;
assign addr[57650]= -1975871368;
assign addr[57651]= -1944661739;
assign addr[57652]= -1910985158;
assign addr[57653]= -1874884346;
assign addr[57654]= -1836405100;
assign addr[57655]= -1795596234;
assign addr[57656]= -1752509516;
assign addr[57657]= -1707199606;
assign addr[57658]= -1659723983;
assign addr[57659]= -1610142873;
assign addr[57660]= -1558519173;
assign addr[57661]= -1504918373;
assign addr[57662]= -1449408469;
assign addr[57663]= -1392059879;
assign addr[57664]= -1332945355;
assign addr[57665]= -1272139887;
assign addr[57666]= -1209720613;
assign addr[57667]= -1145766716;
assign addr[57668]= -1080359326;
assign addr[57669]= -1013581418;
assign addr[57670]= -945517704;
assign addr[57671]= -876254528;
assign addr[57672]= -805879757;
assign addr[57673]= -734482665;
assign addr[57674]= -662153826;
assign addr[57675]= -588984994;
assign addr[57676]= -515068990;
assign addr[57677]= -440499581;
assign addr[57678]= -365371365;
assign addr[57679]= -289779648;
assign addr[57680]= -213820322;
assign addr[57681]= -137589750;
assign addr[57682]= -61184634;
assign addr[57683]= 15298099;
assign addr[57684]= 91761426;
assign addr[57685]= 168108346;
assign addr[57686]= 244242007;
assign addr[57687]= 320065829;
assign addr[57688]= 395483624;
assign addr[57689]= 470399716;
assign addr[57690]= 544719071;
assign addr[57691]= 618347408;
assign addr[57692]= 691191324;
assign addr[57693]= 763158411;
assign addr[57694]= 834157373;
assign addr[57695]= 904098143;
assign addr[57696]= 972891995;
assign addr[57697]= 1040451659;
assign addr[57698]= 1106691431;
assign addr[57699]= 1171527280;
assign addr[57700]= 1234876957;
assign addr[57701]= 1296660098;
assign addr[57702]= 1356798326;
assign addr[57703]= 1415215352;
assign addr[57704]= 1471837070;
assign addr[57705]= 1526591649;
assign addr[57706]= 1579409630;
assign addr[57707]= 1630224009;
assign addr[57708]= 1678970324;
assign addr[57709]= 1725586737;
assign addr[57710]= 1770014111;
assign addr[57711]= 1812196087;
assign addr[57712]= 1852079154;
assign addr[57713]= 1889612716;
assign addr[57714]= 1924749160;
assign addr[57715]= 1957443913;
assign addr[57716]= 1987655498;
assign addr[57717]= 2015345591;
assign addr[57718]= 2040479063;
assign addr[57719]= 2063024031;
assign addr[57720]= 2082951896;
assign addr[57721]= 2100237377;
assign addr[57722]= 2114858546;
assign addr[57723]= 2126796855;
assign addr[57724]= 2136037160;
assign addr[57725]= 2142567738;
assign addr[57726]= 2146380306;
assign addr[57727]= 2147470025;
assign addr[57728]= 2145835515;
assign addr[57729]= 2141478848;
assign addr[57730]= 2134405552;
assign addr[57731]= 2124624598;
assign addr[57732]= 2112148396;
assign addr[57733]= 2096992772;
assign addr[57734]= 2079176953;
assign addr[57735]= 2058723538;
assign addr[57736]= 2035658475;
assign addr[57737]= 2010011024;
assign addr[57738]= 1981813720;
assign addr[57739]= 1951102334;
assign addr[57740]= 1917915825;
assign addr[57741]= 1882296293;
assign addr[57742]= 1844288924;
assign addr[57743]= 1803941934;
assign addr[57744]= 1761306505;
assign addr[57745]= 1716436725;
assign addr[57746]= 1669389513;
assign addr[57747]= 1620224553;
assign addr[57748]= 1569004214;
assign addr[57749]= 1515793473;
assign addr[57750]= 1460659832;
assign addr[57751]= 1403673233;
assign addr[57752]= 1344905966;
assign addr[57753]= 1284432584;
assign addr[57754]= 1222329801;
assign addr[57755]= 1158676398;
assign addr[57756]= 1093553126;
assign addr[57757]= 1027042599;
assign addr[57758]= 959229189;
assign addr[57759]= 890198924;
assign addr[57760]= 820039373;
assign addr[57761]= 748839539;
assign addr[57762]= 676689746;
assign addr[57763]= 603681519;
assign addr[57764]= 529907477;
assign addr[57765]= 455461206;
assign addr[57766]= 380437148;
assign addr[57767]= 304930476;
assign addr[57768]= 229036977;
assign addr[57769]= 152852926;
assign addr[57770]= 76474970;
assign addr[57771]= 0;
assign addr[57772]= -76474970;
assign addr[57773]= -152852926;
assign addr[57774]= -229036977;
assign addr[57775]= -304930476;
assign addr[57776]= -380437148;
assign addr[57777]= -455461206;
assign addr[57778]= -529907477;
assign addr[57779]= -603681519;
assign addr[57780]= -676689746;
assign addr[57781]= -748839539;
assign addr[57782]= -820039373;
assign addr[57783]= -890198924;
assign addr[57784]= -959229189;
assign addr[57785]= -1027042599;
assign addr[57786]= -1093553126;
assign addr[57787]= -1158676398;
assign addr[57788]= -1222329801;
assign addr[57789]= -1284432584;
assign addr[57790]= -1344905966;
assign addr[57791]= -1403673233;
assign addr[57792]= -1460659832;
assign addr[57793]= -1515793473;
assign addr[57794]= -1569004214;
assign addr[57795]= -1620224553;
assign addr[57796]= -1669389513;
assign addr[57797]= -1716436725;
assign addr[57798]= -1761306505;
assign addr[57799]= -1803941934;
assign addr[57800]= -1844288924;
assign addr[57801]= -1882296293;
assign addr[57802]= -1917915825;
assign addr[57803]= -1951102334;
assign addr[57804]= -1981813720;
assign addr[57805]= -2010011024;
assign addr[57806]= -2035658475;
assign addr[57807]= -2058723538;
assign addr[57808]= -2079176953;
assign addr[57809]= -2096992772;
assign addr[57810]= -2112148396;
assign addr[57811]= -2124624598;
assign addr[57812]= -2134405552;
assign addr[57813]= -2141478848;
assign addr[57814]= -2145835515;
assign addr[57815]= -2147470025;
assign addr[57816]= -2146380306;
assign addr[57817]= -2142567738;
assign addr[57818]= -2136037160;
assign addr[57819]= -2126796855;
assign addr[57820]= -2114858546;
assign addr[57821]= -2100237377;
assign addr[57822]= -2082951896;
assign addr[57823]= -2063024031;
assign addr[57824]= -2040479063;
assign addr[57825]= -2015345591;
assign addr[57826]= -1987655498;
assign addr[57827]= -1957443913;
assign addr[57828]= -1924749160;
assign addr[57829]= -1889612716;
assign addr[57830]= -1852079154;
assign addr[57831]= -1812196087;
assign addr[57832]= -1770014111;
assign addr[57833]= -1725586737;
assign addr[57834]= -1678970324;
assign addr[57835]= -1630224009;
assign addr[57836]= -1579409630;
assign addr[57837]= -1526591649;
assign addr[57838]= -1471837070;
assign addr[57839]= -1415215352;
assign addr[57840]= -1356798326;
assign addr[57841]= -1296660098;
assign addr[57842]= -1234876957;
assign addr[57843]= -1171527280;
assign addr[57844]= -1106691431;
assign addr[57845]= -1040451659;
assign addr[57846]= -972891995;
assign addr[57847]= -904098143;
assign addr[57848]= -834157373;
assign addr[57849]= -763158411;
assign addr[57850]= -691191324;
assign addr[57851]= -618347408;
assign addr[57852]= -544719071;
assign addr[57853]= -470399716;
assign addr[57854]= -395483624;
assign addr[57855]= -320065829;
assign addr[57856]= -244242007;
assign addr[57857]= -168108346;
assign addr[57858]= -91761426;
assign addr[57859]= -15298099;
assign addr[57860]= 61184634;
assign addr[57861]= 137589750;
assign addr[57862]= 213820322;
assign addr[57863]= 289779648;
assign addr[57864]= 365371365;
assign addr[57865]= 440499581;
assign addr[57866]= 515068990;
assign addr[57867]= 588984994;
assign addr[57868]= 662153826;
assign addr[57869]= 734482665;
assign addr[57870]= 805879757;
assign addr[57871]= 876254528;
assign addr[57872]= 945517704;
assign addr[57873]= 1013581418;
assign addr[57874]= 1080359326;
assign addr[57875]= 1145766716;
assign addr[57876]= 1209720613;
assign addr[57877]= 1272139887;
assign addr[57878]= 1332945355;
assign addr[57879]= 1392059879;
assign addr[57880]= 1449408469;
assign addr[57881]= 1504918373;
assign addr[57882]= 1558519173;
assign addr[57883]= 1610142873;
assign addr[57884]= 1659723983;
assign addr[57885]= 1707199606;
assign addr[57886]= 1752509516;
assign addr[57887]= 1795596234;
assign addr[57888]= 1836405100;
assign addr[57889]= 1874884346;
assign addr[57890]= 1910985158;
assign addr[57891]= 1944661739;
assign addr[57892]= 1975871368;
assign addr[57893]= 2004574453;
assign addr[57894]= 2030734582;
assign addr[57895]= 2054318569;
assign addr[57896]= 2075296495;
assign addr[57897]= 2093641749;
assign addr[57898]= 2109331059;
assign addr[57899]= 2122344521;
assign addr[57900]= 2132665626;
assign addr[57901]= 2140281282;
assign addr[57902]= 2145181827;
assign addr[57903]= 2147361045;
assign addr[57904]= 2146816171;
assign addr[57905]= 2143547897;
assign addr[57906]= 2137560369;
assign addr[57907]= 2128861181;
assign addr[57908]= 2117461370;
assign addr[57909]= 2103375398;
assign addr[57910]= 2086621133;
assign addr[57911]= 2067219829;
assign addr[57912]= 2045196100;
assign addr[57913]= 2020577882;
assign addr[57914]= 1993396407;
assign addr[57915]= 1963686155;
assign addr[57916]= 1931484818;
assign addr[57917]= 1896833245;
assign addr[57918]= 1859775393;
assign addr[57919]= 1820358275;
assign addr[57920]= 1778631892;
assign addr[57921]= 1734649179;
assign addr[57922]= 1688465931;
assign addr[57923]= 1640140734;
assign addr[57924]= 1589734894;
assign addr[57925]= 1537312353;
assign addr[57926]= 1482939614;
assign addr[57927]= 1426685652;
assign addr[57928]= 1368621831;
assign addr[57929]= 1308821808;
assign addr[57930]= 1247361445;
assign addr[57931]= 1184318708;
assign addr[57932]= 1119773573;
assign addr[57933]= 1053807919;
assign addr[57934]= 986505429;
assign addr[57935]= 917951481;
assign addr[57936]= 848233042;
assign addr[57937]= 777438554;
assign addr[57938]= 705657826;
assign addr[57939]= 632981917;
assign addr[57940]= 559503022;
assign addr[57941]= 485314355;
assign addr[57942]= 410510029;
assign addr[57943]= 335184940;
assign addr[57944]= 259434643;
assign addr[57945]= 183355234;
assign addr[57946]= 107043224;
assign addr[57947]= 30595422;
assign addr[57948]= -45891193;
assign addr[57949]= -122319591;
assign addr[57950]= -198592817;
assign addr[57951]= -274614114;
assign addr[57952]= -350287041;
assign addr[57953]= -425515602;
assign addr[57954]= -500204365;
assign addr[57955]= -574258580;
assign addr[57956]= -647584304;
assign addr[57957]= -720088517;
assign addr[57958]= -791679244;
assign addr[57959]= -862265664;
assign addr[57960]= -931758235;
assign addr[57961]= -1000068799;
assign addr[57962]= -1067110699;
assign addr[57963]= -1132798888;
assign addr[57964]= -1197050035;
assign addr[57965]= -1259782632;
assign addr[57966]= -1320917099;
assign addr[57967]= -1380375881;
assign addr[57968]= -1438083551;
assign addr[57969]= -1493966902;
assign addr[57970]= -1547955041;
assign addr[57971]= -1599979481;
assign addr[57972]= -1649974225;
assign addr[57973]= -1697875851;
assign addr[57974]= -1743623590;
assign addr[57975]= -1787159411;
assign addr[57976]= -1828428082;
assign addr[57977]= -1867377253;
assign addr[57978]= -1903957513;
assign addr[57979]= -1938122457;
assign addr[57980]= -1969828744;
assign addr[57981]= -1999036154;
assign addr[57982]= -2025707632;
assign addr[57983]= -2049809346;
assign addr[57984]= -2071310720;
assign addr[57985]= -2090184478;
assign addr[57986]= -2106406677;
assign addr[57987]= -2119956737;
assign addr[57988]= -2130817471;
assign addr[57989]= -2138975100;
assign addr[57990]= -2144419275;
assign addr[57991]= -2147143090;
assign addr[57992]= -2147143090;
assign addr[57993]= -2144419275;
assign addr[57994]= -2138975100;
assign addr[57995]= -2130817471;
assign addr[57996]= -2119956737;
assign addr[57997]= -2106406677;
assign addr[57998]= -2090184478;
assign addr[57999]= -2071310720;
assign addr[58000]= -2049809346;
assign addr[58001]= -2025707632;
assign addr[58002]= -1999036154;
assign addr[58003]= -1969828744;
assign addr[58004]= -1938122457;
assign addr[58005]= -1903957513;
assign addr[58006]= -1867377253;
assign addr[58007]= -1828428082;
assign addr[58008]= -1787159411;
assign addr[58009]= -1743623590;
assign addr[58010]= -1697875851;
assign addr[58011]= -1649974225;
assign addr[58012]= -1599979481;
assign addr[58013]= -1547955041;
assign addr[58014]= -1493966902;
assign addr[58015]= -1438083551;
assign addr[58016]= -1380375881;
assign addr[58017]= -1320917099;
assign addr[58018]= -1259782632;
assign addr[58019]= -1197050035;
assign addr[58020]= -1132798888;
assign addr[58021]= -1067110699;
assign addr[58022]= -1000068799;
assign addr[58023]= -931758235;
assign addr[58024]= -862265664;
assign addr[58025]= -791679244;
assign addr[58026]= -720088517;
assign addr[58027]= -647584304;
assign addr[58028]= -574258580;
assign addr[58029]= -500204365;
assign addr[58030]= -425515602;
assign addr[58031]= -350287041;
assign addr[58032]= -274614114;
assign addr[58033]= -198592817;
assign addr[58034]= -122319591;
assign addr[58035]= -45891193;
assign addr[58036]= 30595422;
assign addr[58037]= 107043224;
assign addr[58038]= 183355234;
assign addr[58039]= 259434643;
assign addr[58040]= 335184940;
assign addr[58041]= 410510029;
assign addr[58042]= 485314355;
assign addr[58043]= 559503022;
assign addr[58044]= 632981917;
assign addr[58045]= 705657826;
assign addr[58046]= 777438554;
assign addr[58047]= 848233042;
assign addr[58048]= 917951481;
assign addr[58049]= 986505429;
assign addr[58050]= 1053807919;
assign addr[58051]= 1119773573;
assign addr[58052]= 1184318708;
assign addr[58053]= 1247361445;
assign addr[58054]= 1308821808;
assign addr[58055]= 1368621831;
assign addr[58056]= 1426685652;
assign addr[58057]= 1482939614;
assign addr[58058]= 1537312353;
assign addr[58059]= 1589734894;
assign addr[58060]= 1640140734;
assign addr[58061]= 1688465931;
assign addr[58062]= 1734649179;
assign addr[58063]= 1778631892;
assign addr[58064]= 1820358275;
assign addr[58065]= 1859775393;
assign addr[58066]= 1896833245;
assign addr[58067]= 1931484818;
assign addr[58068]= 1963686155;
assign addr[58069]= 1993396407;
assign addr[58070]= 2020577882;
assign addr[58071]= 2045196100;
assign addr[58072]= 2067219829;
assign addr[58073]= 2086621133;
assign addr[58074]= 2103375398;
assign addr[58075]= 2117461370;
assign addr[58076]= 2128861181;
assign addr[58077]= 2137560369;
assign addr[58078]= 2143547897;
assign addr[58079]= 2146816171;
assign addr[58080]= 2147361045;
assign addr[58081]= 2145181827;
assign addr[58082]= 2140281282;
assign addr[58083]= 2132665626;
assign addr[58084]= 2122344521;
assign addr[58085]= 2109331059;
assign addr[58086]= 2093641749;
assign addr[58087]= 2075296495;
assign addr[58088]= 2054318569;
assign addr[58089]= 2030734582;
assign addr[58090]= 2004574453;
assign addr[58091]= 1975871368;
assign addr[58092]= 1944661739;
assign addr[58093]= 1910985158;
assign addr[58094]= 1874884346;
assign addr[58095]= 1836405100;
assign addr[58096]= 1795596234;
assign addr[58097]= 1752509516;
assign addr[58098]= 1707199606;
assign addr[58099]= 1659723983;
assign addr[58100]= 1610142873;
assign addr[58101]= 1558519173;
assign addr[58102]= 1504918373;
assign addr[58103]= 1449408469;
assign addr[58104]= 1392059879;
assign addr[58105]= 1332945355;
assign addr[58106]= 1272139887;
assign addr[58107]= 1209720613;
assign addr[58108]= 1145766716;
assign addr[58109]= 1080359326;
assign addr[58110]= 1013581418;
assign addr[58111]= 945517704;
assign addr[58112]= 876254528;
assign addr[58113]= 805879757;
assign addr[58114]= 734482665;
assign addr[58115]= 662153826;
assign addr[58116]= 588984994;
assign addr[58117]= 515068990;
assign addr[58118]= 440499581;
assign addr[58119]= 365371365;
assign addr[58120]= 289779648;
assign addr[58121]= 213820322;
assign addr[58122]= 137589750;
assign addr[58123]= 61184634;
assign addr[58124]= -15298099;
assign addr[58125]= -91761426;
assign addr[58126]= -168108346;
assign addr[58127]= -244242007;
assign addr[58128]= -320065829;
assign addr[58129]= -395483624;
assign addr[58130]= -470399716;
assign addr[58131]= -544719071;
assign addr[58132]= -618347408;
assign addr[58133]= -691191324;
assign addr[58134]= -763158411;
assign addr[58135]= -834157373;
assign addr[58136]= -904098143;
assign addr[58137]= -972891995;
assign addr[58138]= -1040451659;
assign addr[58139]= -1106691431;
assign addr[58140]= -1171527280;
assign addr[58141]= -1234876957;
assign addr[58142]= -1296660098;
assign addr[58143]= -1356798326;
assign addr[58144]= -1415215352;
assign addr[58145]= -1471837070;
assign addr[58146]= -1526591649;
assign addr[58147]= -1579409630;
assign addr[58148]= -1630224009;
assign addr[58149]= -1678970324;
assign addr[58150]= -1725586737;
assign addr[58151]= -1770014111;
assign addr[58152]= -1812196087;
assign addr[58153]= -1852079154;
assign addr[58154]= -1889612716;
assign addr[58155]= -1924749160;
assign addr[58156]= -1957443913;
assign addr[58157]= -1987655498;
assign addr[58158]= -2015345591;
assign addr[58159]= -2040479063;
assign addr[58160]= -2063024031;
assign addr[58161]= -2082951896;
assign addr[58162]= -2100237377;
assign addr[58163]= -2114858546;
assign addr[58164]= -2126796855;
assign addr[58165]= -2136037160;
assign addr[58166]= -2142567738;
assign addr[58167]= -2146380306;
assign addr[58168]= -2147470025;
assign addr[58169]= -2145835515;
assign addr[58170]= -2141478848;
assign addr[58171]= -2134405552;
assign addr[58172]= -2124624598;
assign addr[58173]= -2112148396;
assign addr[58174]= -2096992772;
assign addr[58175]= -2079176953;
assign addr[58176]= -2058723538;
assign addr[58177]= -2035658475;
assign addr[58178]= -2010011024;
assign addr[58179]= -1981813720;
assign addr[58180]= -1951102334;
assign addr[58181]= -1917915825;
assign addr[58182]= -1882296293;
assign addr[58183]= -1844288924;
assign addr[58184]= -1803941934;
assign addr[58185]= -1761306505;
assign addr[58186]= -1716436725;
assign addr[58187]= -1669389513;
assign addr[58188]= -1620224553;
assign addr[58189]= -1569004214;
assign addr[58190]= -1515793473;
assign addr[58191]= -1460659832;
assign addr[58192]= -1403673233;
assign addr[58193]= -1344905966;
assign addr[58194]= -1284432584;
assign addr[58195]= -1222329801;
assign addr[58196]= -1158676398;
assign addr[58197]= -1093553126;
assign addr[58198]= -1027042599;
assign addr[58199]= -959229189;
assign addr[58200]= -890198924;
assign addr[58201]= -820039373;
assign addr[58202]= -748839539;
assign addr[58203]= -676689746;
assign addr[58204]= -603681519;
assign addr[58205]= -529907477;
assign addr[58206]= -455461206;
assign addr[58207]= -380437148;
assign addr[58208]= -304930476;
assign addr[58209]= -229036977;
assign addr[58210]= -152852926;
assign addr[58211]= -76474970;
assign addr[58212]= 0;
assign addr[58213]= 76474970;
assign addr[58214]= 152852926;
assign addr[58215]= 229036977;
assign addr[58216]= 304930476;
assign addr[58217]= 380437148;
assign addr[58218]= 455461206;
assign addr[58219]= 529907477;
assign addr[58220]= 603681519;
assign addr[58221]= 676689746;
assign addr[58222]= 748839539;
assign addr[58223]= 820039373;
assign addr[58224]= 890198924;
assign addr[58225]= 959229189;
assign addr[58226]= 1027042599;
assign addr[58227]= 1093553126;
assign addr[58228]= 1158676398;
assign addr[58229]= 1222329801;
assign addr[58230]= 1284432584;
assign addr[58231]= 1344905966;
assign addr[58232]= 1403673233;
assign addr[58233]= 1460659832;
assign addr[58234]= 1515793473;
assign addr[58235]= 1569004214;
assign addr[58236]= 1620224553;
assign addr[58237]= 1669389513;
assign addr[58238]= 1716436725;
assign addr[58239]= 1761306505;
assign addr[58240]= 1803941934;
assign addr[58241]= 1844288924;
assign addr[58242]= 1882296293;
assign addr[58243]= 1917915825;
assign addr[58244]= 1951102334;
assign addr[58245]= 1981813720;
assign addr[58246]= 2010011024;
assign addr[58247]= 2035658475;
assign addr[58248]= 2058723538;
assign addr[58249]= 2079176953;
assign addr[58250]= 2096992772;
assign addr[58251]= 2112148396;
assign addr[58252]= 2124624598;
assign addr[58253]= 2134405552;
assign addr[58254]= 2141478848;
assign addr[58255]= 2145835515;
assign addr[58256]= 2147470025;
assign addr[58257]= 2146380306;
assign addr[58258]= 2142567738;
assign addr[58259]= 2136037160;
assign addr[58260]= 2126796855;
assign addr[58261]= 2114858546;
assign addr[58262]= 2100237377;
assign addr[58263]= 2082951896;
assign addr[58264]= 2063024031;
assign addr[58265]= 2040479063;
assign addr[58266]= 2015345591;
assign addr[58267]= 1987655498;
assign addr[58268]= 1957443913;
assign addr[58269]= 1924749160;
assign addr[58270]= 1889612716;
assign addr[58271]= 1852079154;
assign addr[58272]= 1812196087;
assign addr[58273]= 1770014111;
assign addr[58274]= 1725586737;
assign addr[58275]= 1678970324;
assign addr[58276]= 1630224009;
assign addr[58277]= 1579409630;
assign addr[58278]= 1526591649;
assign addr[58279]= 1471837070;
assign addr[58280]= 1415215352;
assign addr[58281]= 1356798326;
assign addr[58282]= 1296660098;
assign addr[58283]= 1234876957;
assign addr[58284]= 1171527280;
assign addr[58285]= 1106691431;
assign addr[58286]= 1040451659;
assign addr[58287]= 972891995;
assign addr[58288]= 904098143;
assign addr[58289]= 834157373;
assign addr[58290]= 763158411;
assign addr[58291]= 691191324;
assign addr[58292]= 618347408;
assign addr[58293]= 544719071;
assign addr[58294]= 470399716;
assign addr[58295]= 395483624;
assign addr[58296]= 320065829;
assign addr[58297]= 244242007;
assign addr[58298]= 168108346;
assign addr[58299]= 91761426;
assign addr[58300]= 15298099;
assign addr[58301]= -61184634;
assign addr[58302]= -137589750;
assign addr[58303]= -213820322;
assign addr[58304]= -289779648;
assign addr[58305]= -365371365;
assign addr[58306]= -440499581;
assign addr[58307]= -515068990;
assign addr[58308]= -588984994;
assign addr[58309]= -662153826;
assign addr[58310]= -734482665;
assign addr[58311]= -805879757;
assign addr[58312]= -876254528;
assign addr[58313]= -945517704;
assign addr[58314]= -1013581418;
assign addr[58315]= -1080359326;
assign addr[58316]= -1145766716;
assign addr[58317]= -1209720613;
assign addr[58318]= -1272139887;
assign addr[58319]= -1332945355;
assign addr[58320]= -1392059879;
assign addr[58321]= -1449408469;
assign addr[58322]= -1504918373;
assign addr[58323]= -1558519173;
assign addr[58324]= -1610142873;
assign addr[58325]= -1659723983;
assign addr[58326]= -1707199606;
assign addr[58327]= -1752509516;
assign addr[58328]= -1795596234;
assign addr[58329]= -1836405100;
assign addr[58330]= -1874884346;
assign addr[58331]= -1910985158;
assign addr[58332]= -1944661739;
assign addr[58333]= -1975871368;
assign addr[58334]= -2004574453;
assign addr[58335]= -2030734582;
assign addr[58336]= -2054318569;
assign addr[58337]= -2075296495;
assign addr[58338]= -2093641749;
assign addr[58339]= -2109331059;
assign addr[58340]= -2122344521;
assign addr[58341]= -2132665626;
assign addr[58342]= -2140281282;
assign addr[58343]= -2145181827;
assign addr[58344]= -2147361045;
assign addr[58345]= -2146816171;
assign addr[58346]= -2143547897;
assign addr[58347]= -2137560369;
assign addr[58348]= -2128861181;
assign addr[58349]= -2117461370;
assign addr[58350]= -2103375398;
assign addr[58351]= -2086621133;
assign addr[58352]= -2067219829;
assign addr[58353]= -2045196100;
assign addr[58354]= -2020577882;
assign addr[58355]= -1993396407;
assign addr[58356]= -1963686155;
assign addr[58357]= -1931484818;
assign addr[58358]= -1896833245;
assign addr[58359]= -1859775393;
assign addr[58360]= -1820358275;
assign addr[58361]= -1778631892;
assign addr[58362]= -1734649179;
assign addr[58363]= -1688465931;
assign addr[58364]= -1640140734;
assign addr[58365]= -1589734894;
assign addr[58366]= -1537312353;
assign addr[58367]= -1482939614;
assign addr[58368]= -1426685652;
assign addr[58369]= -1368621831;
assign addr[58370]= -1308821808;
assign addr[58371]= -1247361445;
assign addr[58372]= -1184318708;
assign addr[58373]= -1119773573;
assign addr[58374]= -1053807919;
assign addr[58375]= -986505429;
assign addr[58376]= -917951481;
assign addr[58377]= -848233042;
assign addr[58378]= -777438554;
assign addr[58379]= -705657826;
assign addr[58380]= -632981917;
assign addr[58381]= -559503022;
assign addr[58382]= -485314355;
assign addr[58383]= -410510029;
assign addr[58384]= -335184940;
assign addr[58385]= -259434643;
assign addr[58386]= -183355234;
assign addr[58387]= -107043224;
assign addr[58388]= -30595422;
assign addr[58389]= 45891193;
assign addr[58390]= 122319591;
assign addr[58391]= 198592817;
assign addr[58392]= 274614114;
assign addr[58393]= 350287041;
assign addr[58394]= 425515602;
assign addr[58395]= 500204365;
assign addr[58396]= 574258580;
assign addr[58397]= 647584304;
assign addr[58398]= 720088517;
assign addr[58399]= 791679244;
assign addr[58400]= 862265664;
assign addr[58401]= 931758235;
assign addr[58402]= 1000068799;
assign addr[58403]= 1067110699;
assign addr[58404]= 1132798888;
assign addr[58405]= 1197050035;
assign addr[58406]= 1259782632;
assign addr[58407]= 1320917099;
assign addr[58408]= 1380375881;
assign addr[58409]= 1438083551;
assign addr[58410]= 1493966902;
assign addr[58411]= 1547955041;
assign addr[58412]= 1599979481;
assign addr[58413]= 1649974225;
assign addr[58414]= 1697875851;
assign addr[58415]= 1743623590;
assign addr[58416]= 1787159411;
assign addr[58417]= 1828428082;
assign addr[58418]= 1867377253;
assign addr[58419]= 1903957513;
assign addr[58420]= 1938122457;
assign addr[58421]= 1969828744;
assign addr[58422]= 1999036154;
assign addr[58423]= 2025707632;
assign addr[58424]= 2049809346;
assign addr[58425]= 2071310720;
assign addr[58426]= 2090184478;
assign addr[58427]= 2106406677;
assign addr[58428]= 2119956737;
assign addr[58429]= 2130817471;
assign addr[58430]= 2138975100;
assign addr[58431]= 2144419275;
assign addr[58432]= 2147143090;
assign addr[58433]= 2147143090;
assign addr[58434]= 2144419275;
assign addr[58435]= 2138975100;
assign addr[58436]= 2130817471;
assign addr[58437]= 2119956737;
assign addr[58438]= 2106406677;
assign addr[58439]= 2090184478;
assign addr[58440]= 2071310720;
assign addr[58441]= 2049809346;
assign addr[58442]= 2025707632;
assign addr[58443]= 1999036154;
assign addr[58444]= 1969828744;
assign addr[58445]= 1938122457;
assign addr[58446]= 1903957513;
assign addr[58447]= 1867377253;
assign addr[58448]= 1828428082;
assign addr[58449]= 1787159411;
assign addr[58450]= 1743623590;
assign addr[58451]= 1697875851;
assign addr[58452]= 1649974225;
assign addr[58453]= 1599979481;
assign addr[58454]= 1547955041;
assign addr[58455]= 1493966902;
assign addr[58456]= 1438083551;
assign addr[58457]= 1380375881;
assign addr[58458]= 1320917099;
assign addr[58459]= 1259782632;
assign addr[58460]= 1197050035;
assign addr[58461]= 1132798888;
assign addr[58462]= 1067110699;
assign addr[58463]= 1000068799;
assign addr[58464]= 931758235;
assign addr[58465]= 862265664;
assign addr[58466]= 791679244;
assign addr[58467]= 720088517;
assign addr[58468]= 647584304;
assign addr[58469]= 574258580;
assign addr[58470]= 500204365;
assign addr[58471]= 425515602;
assign addr[58472]= 350287041;
assign addr[58473]= 274614114;
assign addr[58474]= 198592817;
assign addr[58475]= 122319591;
assign addr[58476]= 45891193;
assign addr[58477]= -30595422;
assign addr[58478]= -107043224;
assign addr[58479]= -183355234;
assign addr[58480]= -259434643;
assign addr[58481]= -335184940;
assign addr[58482]= -410510029;
assign addr[58483]= -485314355;
assign addr[58484]= -559503022;
assign addr[58485]= -632981917;
assign addr[58486]= -705657826;
assign addr[58487]= -777438554;
assign addr[58488]= -848233042;
assign addr[58489]= -917951481;
assign addr[58490]= -986505429;
assign addr[58491]= -1053807919;
assign addr[58492]= -1119773573;
assign addr[58493]= -1184318708;
assign addr[58494]= -1247361445;
assign addr[58495]= -1308821808;
assign addr[58496]= -1368621831;
assign addr[58497]= -1426685652;
assign addr[58498]= -1482939614;
assign addr[58499]= -1537312353;
assign addr[58500]= -1589734894;
assign addr[58501]= -1640140734;
assign addr[58502]= -1688465931;
assign addr[58503]= -1734649179;
assign addr[58504]= -1778631892;
assign addr[58505]= -1820358275;
assign addr[58506]= -1859775393;
assign addr[58507]= -1896833245;
assign addr[58508]= -1931484818;
assign addr[58509]= -1963686155;
assign addr[58510]= -1993396407;
assign addr[58511]= -2020577882;
assign addr[58512]= -2045196100;
assign addr[58513]= -2067219829;
assign addr[58514]= -2086621133;
assign addr[58515]= -2103375398;
assign addr[58516]= -2117461370;
assign addr[58517]= -2128861181;
assign addr[58518]= -2137560369;
assign addr[58519]= -2143547897;
assign addr[58520]= -2146816171;
assign addr[58521]= -2147361045;
assign addr[58522]= -2145181827;
assign addr[58523]= -2140281282;
assign addr[58524]= -2132665626;
assign addr[58525]= -2122344521;
assign addr[58526]= -2109331059;
assign addr[58527]= -2093641749;
assign addr[58528]= -2075296495;
assign addr[58529]= -2054318569;
assign addr[58530]= -2030734582;
assign addr[58531]= -2004574453;
assign addr[58532]= -1975871368;
assign addr[58533]= -1944661739;
assign addr[58534]= -1910985158;
assign addr[58535]= -1874884346;
assign addr[58536]= -1836405100;
assign addr[58537]= -1795596234;
assign addr[58538]= -1752509516;
assign addr[58539]= -1707199606;
assign addr[58540]= -1659723983;
assign addr[58541]= -1610142873;
assign addr[58542]= -1558519173;
assign addr[58543]= -1504918373;
assign addr[58544]= -1449408469;
assign addr[58545]= -1392059879;
assign addr[58546]= -1332945355;
assign addr[58547]= -1272139887;
assign addr[58548]= -1209720613;
assign addr[58549]= -1145766716;
assign addr[58550]= -1080359326;
assign addr[58551]= -1013581418;
assign addr[58552]= -945517704;
assign addr[58553]= -876254528;
assign addr[58554]= -805879757;
assign addr[58555]= -734482665;
assign addr[58556]= -662153826;
assign addr[58557]= -588984994;
assign addr[58558]= -515068990;
assign addr[58559]= -440499581;
assign addr[58560]= -365371365;
assign addr[58561]= -289779648;
assign addr[58562]= -213820322;
assign addr[58563]= -137589750;
assign addr[58564]= -61184634;
assign addr[58565]= 15298099;
assign addr[58566]= 91761426;
assign addr[58567]= 168108346;
assign addr[58568]= 244242007;
assign addr[58569]= 320065829;
assign addr[58570]= 395483624;
assign addr[58571]= 470399716;
assign addr[58572]= 544719071;
assign addr[58573]= 618347408;
assign addr[58574]= 691191324;
assign addr[58575]= 763158411;
assign addr[58576]= 834157373;
assign addr[58577]= 904098143;
assign addr[58578]= 972891995;
assign addr[58579]= 1040451659;
assign addr[58580]= 1106691431;
assign addr[58581]= 1171527280;
assign addr[58582]= 1234876957;
assign addr[58583]= 1296660098;
assign addr[58584]= 1356798326;
assign addr[58585]= 1415215352;
assign addr[58586]= 1471837070;
assign addr[58587]= 1526591649;
assign addr[58588]= 1579409630;
assign addr[58589]= 1630224009;
assign addr[58590]= 1678970324;
assign addr[58591]= 1725586737;
assign addr[58592]= 1770014111;
assign addr[58593]= 1812196087;
assign addr[58594]= 1852079154;
assign addr[58595]= 1889612716;
assign addr[58596]= 1924749160;
assign addr[58597]= 1957443913;
assign addr[58598]= 1987655498;
assign addr[58599]= 2015345591;
assign addr[58600]= 2040479063;
assign addr[58601]= 2063024031;
assign addr[58602]= 2082951896;
assign addr[58603]= 2100237377;
assign addr[58604]= 2114858546;
assign addr[58605]= 2126796855;
assign addr[58606]= 2136037160;
assign addr[58607]= 2142567738;
assign addr[58608]= 2146380306;
assign addr[58609]= 2147470025;
assign addr[58610]= 2145835515;
assign addr[58611]= 2141478848;
assign addr[58612]= 2134405552;
assign addr[58613]= 2124624598;
assign addr[58614]= 2112148396;
assign addr[58615]= 2096992772;
assign addr[58616]= 2079176953;
assign addr[58617]= 2058723538;
assign addr[58618]= 2035658475;
assign addr[58619]= 2010011024;
assign addr[58620]= 1981813720;
assign addr[58621]= 1951102334;
assign addr[58622]= 1917915825;
assign addr[58623]= 1882296293;
assign addr[58624]= 1844288924;
assign addr[58625]= 1803941934;
assign addr[58626]= 1761306505;
assign addr[58627]= 1716436725;
assign addr[58628]= 1669389513;
assign addr[58629]= 1620224553;
assign addr[58630]= 1569004214;
assign addr[58631]= 1515793473;
assign addr[58632]= 1460659832;
assign addr[58633]= 1403673233;
assign addr[58634]= 1344905966;
assign addr[58635]= 1284432584;
assign addr[58636]= 1222329801;
assign addr[58637]= 1158676398;
assign addr[58638]= 1093553126;
assign addr[58639]= 1027042599;
assign addr[58640]= 959229189;
assign addr[58641]= 890198924;
assign addr[58642]= 820039373;
assign addr[58643]= 748839539;
assign addr[58644]= 676689746;
assign addr[58645]= 603681519;
assign addr[58646]= 529907477;
assign addr[58647]= 455461206;
assign addr[58648]= 380437148;
assign addr[58649]= 304930476;
assign addr[58650]= 229036977;
assign addr[58651]= 152852926;
assign addr[58652]= 76474970;
assign addr[58653]= 0;
assign addr[58654]= -76474970;
assign addr[58655]= -152852926;
assign addr[58656]= -229036977;
assign addr[58657]= -304930476;
assign addr[58658]= -380437148;
assign addr[58659]= -455461206;
assign addr[58660]= -529907477;
assign addr[58661]= -603681519;
assign addr[58662]= -676689746;
assign addr[58663]= -748839539;
assign addr[58664]= -820039373;
assign addr[58665]= -890198924;
assign addr[58666]= -959229189;
assign addr[58667]= -1027042599;
assign addr[58668]= -1093553126;
assign addr[58669]= -1158676398;
assign addr[58670]= -1222329801;
assign addr[58671]= -1284432584;
assign addr[58672]= -1344905966;
assign addr[58673]= -1403673233;
assign addr[58674]= -1460659832;
assign addr[58675]= -1515793473;
assign addr[58676]= -1569004214;
assign addr[58677]= -1620224553;
assign addr[58678]= -1669389513;
assign addr[58679]= -1716436725;
assign addr[58680]= -1761306505;
assign addr[58681]= -1803941934;
assign addr[58682]= -1844288924;
assign addr[58683]= -1882296293;
assign addr[58684]= -1917915825;
assign addr[58685]= -1951102334;
assign addr[58686]= -1981813720;
assign addr[58687]= -2010011024;
assign addr[58688]= -2035658475;
assign addr[58689]= -2058723538;
assign addr[58690]= -2079176953;
assign addr[58691]= -2096992772;
assign addr[58692]= -2112148396;
assign addr[58693]= -2124624598;
assign addr[58694]= -2134405552;
assign addr[58695]= -2141478848;
assign addr[58696]= -2145835515;
assign addr[58697]= -2147470025;
assign addr[58698]= -2146380306;
assign addr[58699]= -2142567738;
assign addr[58700]= -2136037160;
assign addr[58701]= -2126796855;
assign addr[58702]= -2114858546;
assign addr[58703]= -2100237377;
assign addr[58704]= -2082951896;
assign addr[58705]= -2063024031;
assign addr[58706]= -2040479063;
assign addr[58707]= -2015345591;
assign addr[58708]= -1987655498;
assign addr[58709]= -1957443913;
assign addr[58710]= -1924749160;
assign addr[58711]= -1889612716;
assign addr[58712]= -1852079154;
assign addr[58713]= -1812196087;
assign addr[58714]= -1770014111;
assign addr[58715]= -1725586737;
assign addr[58716]= -1678970324;
assign addr[58717]= -1630224009;
assign addr[58718]= -1579409630;
assign addr[58719]= -1526591649;
assign addr[58720]= -1471837070;
assign addr[58721]= -1415215352;
assign addr[58722]= -1356798326;
assign addr[58723]= -1296660098;
assign addr[58724]= -1234876957;
assign addr[58725]= -1171527280;
assign addr[58726]= -1106691431;
assign addr[58727]= -1040451659;
assign addr[58728]= -972891995;
assign addr[58729]= -904098143;
assign addr[58730]= -834157373;
assign addr[58731]= -763158411;
assign addr[58732]= -691191324;
assign addr[58733]= -618347408;
assign addr[58734]= -544719071;
assign addr[58735]= -470399716;
assign addr[58736]= -395483624;
assign addr[58737]= -320065829;
assign addr[58738]= -244242007;
assign addr[58739]= -168108346;
assign addr[58740]= -91761426;
assign addr[58741]= -15298099;
assign addr[58742]= 61184634;
assign addr[58743]= 137589750;
assign addr[58744]= 213820322;
assign addr[58745]= 289779648;
assign addr[58746]= 365371365;
assign addr[58747]= 440499581;
assign addr[58748]= 515068990;
assign addr[58749]= 588984994;
assign addr[58750]= 662153826;
assign addr[58751]= 734482665;
assign addr[58752]= 805879757;
assign addr[58753]= 876254528;
assign addr[58754]= 945517704;
assign addr[58755]= 1013581418;
assign addr[58756]= 1080359326;
assign addr[58757]= 1145766716;
assign addr[58758]= 1209720613;
assign addr[58759]= 1272139887;
assign addr[58760]= 1332945355;
assign addr[58761]= 1392059879;
assign addr[58762]= 1449408469;
assign addr[58763]= 1504918373;
assign addr[58764]= 1558519173;
assign addr[58765]= 1610142873;
assign addr[58766]= 1659723983;
assign addr[58767]= 1707199606;
assign addr[58768]= 1752509516;
assign addr[58769]= 1795596234;
assign addr[58770]= 1836405100;
assign addr[58771]= 1874884346;
assign addr[58772]= 1910985158;
assign addr[58773]= 1944661739;
assign addr[58774]= 1975871368;
assign addr[58775]= 2004574453;
assign addr[58776]= 2030734582;
assign addr[58777]= 2054318569;
assign addr[58778]= 2075296495;
assign addr[58779]= 2093641749;
assign addr[58780]= 2109331059;
assign addr[58781]= 2122344521;
assign addr[58782]= 2132665626;
assign addr[58783]= 2140281282;
assign addr[58784]= 2145181827;
assign addr[58785]= 2147361045;
assign addr[58786]= 2146816171;
assign addr[58787]= 2143547897;
assign addr[58788]= 2137560369;
assign addr[58789]= 2128861181;
assign addr[58790]= 2117461370;
assign addr[58791]= 2103375398;
assign addr[58792]= 2086621133;
assign addr[58793]= 2067219829;
assign addr[58794]= 2045196100;
assign addr[58795]= 2020577882;
assign addr[58796]= 1993396407;
assign addr[58797]= 1963686155;
assign addr[58798]= 1931484818;
assign addr[58799]= 1896833245;
assign addr[58800]= 1859775393;
assign addr[58801]= 1820358275;
assign addr[58802]= 1778631892;
assign addr[58803]= 1734649179;
assign addr[58804]= 1688465931;
assign addr[58805]= 1640140734;
assign addr[58806]= 1589734894;
assign addr[58807]= 1537312353;
assign addr[58808]= 1482939614;
assign addr[58809]= 1426685652;
assign addr[58810]= 1368621831;
assign addr[58811]= 1308821808;
assign addr[58812]= 1247361445;
assign addr[58813]= 1184318708;
assign addr[58814]= 1119773573;
assign addr[58815]= 1053807919;
assign addr[58816]= 986505429;
assign addr[58817]= 917951481;
assign addr[58818]= 848233042;
assign addr[58819]= 777438554;
assign addr[58820]= 705657826;
assign addr[58821]= 632981917;
assign addr[58822]= 559503022;
assign addr[58823]= 485314355;
assign addr[58824]= 410510029;
assign addr[58825]= 335184940;
assign addr[58826]= 259434643;
assign addr[58827]= 183355234;
assign addr[58828]= 107043224;
assign addr[58829]= 30595422;
assign addr[58830]= -45891193;
assign addr[58831]= -122319591;
assign addr[58832]= -198592817;
assign addr[58833]= -274614114;
assign addr[58834]= -350287041;
assign addr[58835]= -425515602;
assign addr[58836]= -500204365;
assign addr[58837]= -574258580;
assign addr[58838]= -647584304;
assign addr[58839]= -720088517;
assign addr[58840]= -791679244;
assign addr[58841]= -862265664;
assign addr[58842]= -931758235;
assign addr[58843]= -1000068799;
assign addr[58844]= -1067110699;
assign addr[58845]= -1132798888;
assign addr[58846]= -1197050035;
assign addr[58847]= -1259782632;
assign addr[58848]= -1320917099;
assign addr[58849]= -1380375881;
assign addr[58850]= -1438083551;
assign addr[58851]= -1493966902;
assign addr[58852]= -1547955041;
assign addr[58853]= -1599979481;
assign addr[58854]= -1649974225;
assign addr[58855]= -1697875851;
assign addr[58856]= -1743623590;
assign addr[58857]= -1787159411;
assign addr[58858]= -1828428082;
assign addr[58859]= -1867377253;
assign addr[58860]= -1903957513;
assign addr[58861]= -1938122457;
assign addr[58862]= -1969828744;
assign addr[58863]= -1999036154;
assign addr[58864]= -2025707632;
assign addr[58865]= -2049809346;
assign addr[58866]= -2071310720;
assign addr[58867]= -2090184478;
assign addr[58868]= -2106406677;
assign addr[58869]= -2119956737;
assign addr[58870]= -2130817471;
assign addr[58871]= -2138975100;
assign addr[58872]= -2144419275;
assign addr[58873]= -2147143090;
assign addr[58874]= -2147143090;
assign addr[58875]= -2144419275;
assign addr[58876]= -2138975100;
assign addr[58877]= -2130817471;
assign addr[58878]= -2119956737;
assign addr[58879]= -2106406677;
assign addr[58880]= -2090184478;
assign addr[58881]= -2071310720;
assign addr[58882]= -2049809346;
assign addr[58883]= -2025707632;
assign addr[58884]= -1999036154;
assign addr[58885]= -1969828744;
assign addr[58886]= -1938122457;
assign addr[58887]= -1903957513;
assign addr[58888]= -1867377253;
assign addr[58889]= -1828428082;
assign addr[58890]= -1787159411;
assign addr[58891]= -1743623590;
assign addr[58892]= -1697875851;
assign addr[58893]= -1649974225;
assign addr[58894]= -1599979481;
assign addr[58895]= -1547955041;
assign addr[58896]= -1493966902;
assign addr[58897]= -1438083551;
assign addr[58898]= -1380375881;
assign addr[58899]= -1320917099;
assign addr[58900]= -1259782632;
assign addr[58901]= -1197050035;
assign addr[58902]= -1132798888;
assign addr[58903]= -1067110699;
assign addr[58904]= -1000068799;
assign addr[58905]= -931758235;
assign addr[58906]= -862265664;
assign addr[58907]= -791679244;
assign addr[58908]= -720088517;
assign addr[58909]= -647584304;
assign addr[58910]= -574258580;
assign addr[58911]= -500204365;
assign addr[58912]= -425515602;
assign addr[58913]= -350287041;
assign addr[58914]= -274614114;
assign addr[58915]= -198592817;
assign addr[58916]= -122319591;
assign addr[58917]= -45891193;
assign addr[58918]= 30595422;
assign addr[58919]= 107043224;
assign addr[58920]= 183355234;
assign addr[58921]= 259434643;
assign addr[58922]= 335184940;
assign addr[58923]= 410510029;
assign addr[58924]= 485314355;
assign addr[58925]= 559503022;
assign addr[58926]= 632981917;
assign addr[58927]= 705657826;
assign addr[58928]= 777438554;
assign addr[58929]= 848233042;
assign addr[58930]= 917951481;
assign addr[58931]= 986505429;
assign addr[58932]= 1053807919;
assign addr[58933]= 1119773573;
assign addr[58934]= 1184318708;
assign addr[58935]= 1247361445;
assign addr[58936]= 1308821808;
assign addr[58937]= 1368621831;
assign addr[58938]= 1426685652;
assign addr[58939]= 1482939614;
assign addr[58940]= 1537312353;
assign addr[58941]= 1589734894;
assign addr[58942]= 1640140734;
assign addr[58943]= 1688465931;
assign addr[58944]= 1734649179;
assign addr[58945]= 1778631892;
assign addr[58946]= 1820358275;
assign addr[58947]= 1859775393;
assign addr[58948]= 1896833245;
assign addr[58949]= 1931484818;
assign addr[58950]= 1963686155;
assign addr[58951]= 1993396407;
assign addr[58952]= 2020577882;
assign addr[58953]= 2045196100;
assign addr[58954]= 2067219829;
assign addr[58955]= 2086621133;
assign addr[58956]= 2103375398;
assign addr[58957]= 2117461370;
assign addr[58958]= 2128861181;
assign addr[58959]= 2137560369;
assign addr[58960]= 2143547897;
assign addr[58961]= 2146816171;
assign addr[58962]= 2147361045;
assign addr[58963]= 2145181827;
assign addr[58964]= 2140281282;
assign addr[58965]= 2132665626;
assign addr[58966]= 2122344521;
assign addr[58967]= 2109331059;
assign addr[58968]= 2093641749;
assign addr[58969]= 2075296495;
assign addr[58970]= 2054318569;
assign addr[58971]= 2030734582;
assign addr[58972]= 2004574453;
assign addr[58973]= 1975871368;
assign addr[58974]= 1944661739;
assign addr[58975]= 1910985158;
assign addr[58976]= 1874884346;
assign addr[58977]= 1836405100;
assign addr[58978]= 1795596234;
assign addr[58979]= 1752509516;
assign addr[58980]= 1707199606;
assign addr[58981]= 1659723983;
assign addr[58982]= 1610142873;
assign addr[58983]= 1558519173;
assign addr[58984]= 1504918373;
assign addr[58985]= 1449408469;
assign addr[58986]= 1392059879;
assign addr[58987]= 1332945355;
assign addr[58988]= 1272139887;
assign addr[58989]= 1209720613;
assign addr[58990]= 1145766716;
assign addr[58991]= 1080359326;
assign addr[58992]= 1013581418;
assign addr[58993]= 945517704;
assign addr[58994]= 876254528;
assign addr[58995]= 805879757;
assign addr[58996]= 734482665;
assign addr[58997]= 662153826;
assign addr[58998]= 588984994;
assign addr[58999]= 515068990;
assign addr[59000]= 440499581;
assign addr[59001]= 365371365;
assign addr[59002]= 289779648;
assign addr[59003]= 213820322;
assign addr[59004]= 137589750;
assign addr[59005]= 61184634;
assign addr[59006]= -15298099;
assign addr[59007]= -91761426;
assign addr[59008]= -168108346;
assign addr[59009]= -244242007;
assign addr[59010]= -320065829;
assign addr[59011]= -395483624;
assign addr[59012]= -470399716;
assign addr[59013]= -544719071;
assign addr[59014]= -618347408;
assign addr[59015]= -691191324;
assign addr[59016]= -763158411;
assign addr[59017]= -834157373;
assign addr[59018]= -904098143;
assign addr[59019]= -972891995;
assign addr[59020]= -1040451659;
assign addr[59021]= -1106691431;
assign addr[59022]= -1171527280;
assign addr[59023]= -1234876957;
assign addr[59024]= -1296660098;
assign addr[59025]= -1356798326;
assign addr[59026]= -1415215352;
assign addr[59027]= -1471837070;
assign addr[59028]= -1526591649;
assign addr[59029]= -1579409630;
assign addr[59030]= -1630224009;
assign addr[59031]= -1678970324;
assign addr[59032]= -1725586737;
assign addr[59033]= -1770014111;
assign addr[59034]= -1812196087;
assign addr[59035]= -1852079154;
assign addr[59036]= -1889612716;
assign addr[59037]= -1924749160;
assign addr[59038]= -1957443913;
assign addr[59039]= -1987655498;
assign addr[59040]= -2015345591;
assign addr[59041]= -2040479063;
assign addr[59042]= -2063024031;
assign addr[59043]= -2082951896;
assign addr[59044]= -2100237377;
assign addr[59045]= -2114858546;
assign addr[59046]= -2126796855;
assign addr[59047]= -2136037160;
assign addr[59048]= -2142567738;
assign addr[59049]= -2146380306;
assign addr[59050]= -2147470025;
assign addr[59051]= -2145835515;
assign addr[59052]= -2141478848;
assign addr[59053]= -2134405552;
assign addr[59054]= -2124624598;
assign addr[59055]= -2112148396;
assign addr[59056]= -2096992772;
assign addr[59057]= -2079176953;
assign addr[59058]= -2058723538;
assign addr[59059]= -2035658475;
assign addr[59060]= -2010011024;
assign addr[59061]= -1981813720;
assign addr[59062]= -1951102334;
assign addr[59063]= -1917915825;
assign addr[59064]= -1882296293;
assign addr[59065]= -1844288924;
assign addr[59066]= -1803941934;
assign addr[59067]= -1761306505;
assign addr[59068]= -1716436725;
assign addr[59069]= -1669389513;
assign addr[59070]= -1620224553;
assign addr[59071]= -1569004214;
assign addr[59072]= -1515793473;
assign addr[59073]= -1460659832;
assign addr[59074]= -1403673233;
assign addr[59075]= -1344905966;
assign addr[59076]= -1284432584;
assign addr[59077]= -1222329801;
assign addr[59078]= -1158676398;
assign addr[59079]= -1093553126;
assign addr[59080]= -1027042599;
assign addr[59081]= -959229189;
assign addr[59082]= -890198924;
assign addr[59083]= -820039373;
assign addr[59084]= -748839539;
assign addr[59085]= -676689746;
assign addr[59086]= -603681519;
assign addr[59087]= -529907477;
assign addr[59088]= -455461206;
assign addr[59089]= -380437148;
assign addr[59090]= -304930476;
assign addr[59091]= -229036977;
assign addr[59092]= -152852926;
assign addr[59093]= -76474970;
assign addr[59094]= 0;
assign addr[59095]= 76474970;
assign addr[59096]= 152852926;
assign addr[59097]= 229036977;
assign addr[59098]= 304930476;
assign addr[59099]= 380437148;
assign addr[59100]= 455461206;
assign addr[59101]= 529907477;
assign addr[59102]= 603681519;
assign addr[59103]= 676689746;
assign addr[59104]= 748839539;
assign addr[59105]= 820039373;
assign addr[59106]= 890198924;
assign addr[59107]= 959229189;
assign addr[59108]= 1027042599;
assign addr[59109]= 1093553126;
assign addr[59110]= 1158676398;
assign addr[59111]= 1222329801;
assign addr[59112]= 1284432584;
assign addr[59113]= 1344905966;
assign addr[59114]= 1403673233;
assign addr[59115]= 1460659832;
assign addr[59116]= 1515793473;
assign addr[59117]= 1569004214;
assign addr[59118]= 1620224553;
assign addr[59119]= 1669389513;
assign addr[59120]= 1716436725;
assign addr[59121]= 1761306505;
assign addr[59122]= 1803941934;
assign addr[59123]= 1844288924;
assign addr[59124]= 1882296293;
assign addr[59125]= 1917915825;
assign addr[59126]= 1951102334;
assign addr[59127]= 1981813720;
assign addr[59128]= 2010011024;
assign addr[59129]= 2035658475;
assign addr[59130]= 2058723538;
assign addr[59131]= 2079176953;
assign addr[59132]= 2096992772;
assign addr[59133]= 2112148396;
assign addr[59134]= 2124624598;
assign addr[59135]= 2134405552;
assign addr[59136]= 2141478848;
assign addr[59137]= 2145835515;
assign addr[59138]= 2147470025;
assign addr[59139]= 2146380306;
assign addr[59140]= 2142567738;
assign addr[59141]= 2136037160;
assign addr[59142]= 2126796855;
assign addr[59143]= 2114858546;
assign addr[59144]= 2100237377;
assign addr[59145]= 2082951896;
assign addr[59146]= 2063024031;
assign addr[59147]= 2040479063;
assign addr[59148]= 2015345591;
assign addr[59149]= 1987655498;
assign addr[59150]= 1957443913;
assign addr[59151]= 1924749160;
assign addr[59152]= 1889612716;
assign addr[59153]= 1852079154;
assign addr[59154]= 1812196087;
assign addr[59155]= 1770014111;
assign addr[59156]= 1725586737;
assign addr[59157]= 1678970324;
assign addr[59158]= 1630224009;
assign addr[59159]= 1579409630;
assign addr[59160]= 1526591649;
assign addr[59161]= 1471837070;
assign addr[59162]= 1415215352;
assign addr[59163]= 1356798326;
assign addr[59164]= 1296660098;
assign addr[59165]= 1234876957;
assign addr[59166]= 1171527280;
assign addr[59167]= 1106691431;
assign addr[59168]= 1040451659;
assign addr[59169]= 972891995;
assign addr[59170]= 904098143;
assign addr[59171]= 834157373;
assign addr[59172]= 763158411;
assign addr[59173]= 691191324;
assign addr[59174]= 618347408;
assign addr[59175]= 544719071;
assign addr[59176]= 470399716;
assign addr[59177]= 395483624;
assign addr[59178]= 320065829;
assign addr[59179]= 244242007;
assign addr[59180]= 168108346;
assign addr[59181]= 91761426;
assign addr[59182]= 15298099;
assign addr[59183]= -61184634;
assign addr[59184]= -137589750;
assign addr[59185]= -213820322;
assign addr[59186]= -289779648;
assign addr[59187]= -365371365;
assign addr[59188]= -440499581;
assign addr[59189]= -515068990;
assign addr[59190]= -588984994;
assign addr[59191]= -662153826;
assign addr[59192]= -734482665;
assign addr[59193]= -805879757;
assign addr[59194]= -876254528;
assign addr[59195]= -945517704;
assign addr[59196]= -1013581418;
assign addr[59197]= -1080359326;
assign addr[59198]= -1145766716;
assign addr[59199]= -1209720613;
assign addr[59200]= -1272139887;
assign addr[59201]= -1332945355;
assign addr[59202]= -1392059879;
assign addr[59203]= -1449408469;
assign addr[59204]= -1504918373;
assign addr[59205]= -1558519173;
assign addr[59206]= -1610142873;
assign addr[59207]= -1659723983;
assign addr[59208]= -1707199606;
assign addr[59209]= -1752509516;
assign addr[59210]= -1795596234;
assign addr[59211]= -1836405100;
assign addr[59212]= -1874884346;
assign addr[59213]= -1910985158;
assign addr[59214]= -1944661739;
assign addr[59215]= -1975871368;
assign addr[59216]= -2004574453;
assign addr[59217]= -2030734582;
assign addr[59218]= -2054318569;
assign addr[59219]= -2075296495;
assign addr[59220]= -2093641749;
assign addr[59221]= -2109331059;
assign addr[59222]= -2122344521;
assign addr[59223]= -2132665626;
assign addr[59224]= -2140281282;
assign addr[59225]= -2145181827;
assign addr[59226]= -2147361045;
assign addr[59227]= -2146816171;
assign addr[59228]= -2143547897;
assign addr[59229]= -2137560369;
assign addr[59230]= -2128861181;
assign addr[59231]= -2117461370;
assign addr[59232]= -2103375398;
assign addr[59233]= -2086621133;
assign addr[59234]= -2067219829;
assign addr[59235]= -2045196100;
assign addr[59236]= -2020577882;
assign addr[59237]= -1993396407;
assign addr[59238]= -1963686155;
assign addr[59239]= -1931484818;
assign addr[59240]= -1896833245;
assign addr[59241]= -1859775393;
assign addr[59242]= -1820358275;
assign addr[59243]= -1778631892;
assign addr[59244]= -1734649179;
assign addr[59245]= -1688465931;
assign addr[59246]= -1640140734;
assign addr[59247]= -1589734894;
assign addr[59248]= -1537312353;
assign addr[59249]= -1482939614;
assign addr[59250]= -1426685652;
assign addr[59251]= -1368621831;
assign addr[59252]= -1308821808;
assign addr[59253]= -1247361445;
assign addr[59254]= -1184318708;
assign addr[59255]= -1119773573;
assign addr[59256]= -1053807919;
assign addr[59257]= -986505429;
assign addr[59258]= -917951481;
assign addr[59259]= -848233042;
assign addr[59260]= -777438554;
assign addr[59261]= -705657826;
assign addr[59262]= -632981917;
assign addr[59263]= -559503022;
assign addr[59264]= -485314355;
assign addr[59265]= -410510029;
assign addr[59266]= -335184940;
assign addr[59267]= -259434643;
assign addr[59268]= -183355234;
assign addr[59269]= -107043224;
assign addr[59270]= -30595422;
assign addr[59271]= 45891193;
assign addr[59272]= 122319591;
assign addr[59273]= 198592817;
assign addr[59274]= 274614114;
assign addr[59275]= 350287041;
assign addr[59276]= 425515602;
assign addr[59277]= 500204365;
assign addr[59278]= 574258580;
assign addr[59279]= 647584304;
assign addr[59280]= 720088517;
assign addr[59281]= 791679244;
assign addr[59282]= 862265664;
assign addr[59283]= 931758235;
assign addr[59284]= 1000068799;
assign addr[59285]= 1067110699;
assign addr[59286]= 1132798888;
assign addr[59287]= 1197050035;
assign addr[59288]= 1259782632;
assign addr[59289]= 1320917099;
assign addr[59290]= 1380375881;
assign addr[59291]= 1438083551;
assign addr[59292]= 1493966902;
assign addr[59293]= 1547955041;
assign addr[59294]= 1599979481;
assign addr[59295]= 1649974225;
assign addr[59296]= 1697875851;
assign addr[59297]= 1743623590;
assign addr[59298]= 1787159411;
assign addr[59299]= 1828428082;
assign addr[59300]= 1867377253;
assign addr[59301]= 1903957513;
assign addr[59302]= 1938122457;
assign addr[59303]= 1969828744;
assign addr[59304]= 1999036154;
assign addr[59305]= 2025707632;
assign addr[59306]= 2049809346;
assign addr[59307]= 2071310720;
assign addr[59308]= 2090184478;
assign addr[59309]= 2106406677;
assign addr[59310]= 2119956737;
assign addr[59311]= 2130817471;
assign addr[59312]= 2138975100;
assign addr[59313]= 2144419275;
assign addr[59314]= 2147143090;
assign addr[59315]= 2147143090;
assign addr[59316]= 2144419275;
assign addr[59317]= 2138975100;
assign addr[59318]= 2130817471;
assign addr[59319]= 2119956737;
assign addr[59320]= 2106406677;
assign addr[59321]= 2090184478;
assign addr[59322]= 2071310720;
assign addr[59323]= 2049809346;
assign addr[59324]= 2025707632;
assign addr[59325]= 1999036154;
assign addr[59326]= 1969828744;
assign addr[59327]= 1938122457;
assign addr[59328]= 1903957513;
assign addr[59329]= 1867377253;
assign addr[59330]= 1828428082;
assign addr[59331]= 1787159411;
assign addr[59332]= 1743623590;
assign addr[59333]= 1697875851;
assign addr[59334]= 1649974225;
assign addr[59335]= 1599979481;
assign addr[59336]= 1547955041;
assign addr[59337]= 1493966902;
assign addr[59338]= 1438083551;
assign addr[59339]= 1380375881;
assign addr[59340]= 1320917099;
assign addr[59341]= 1259782632;
assign addr[59342]= 1197050035;
assign addr[59343]= 1132798888;
assign addr[59344]= 1067110699;
assign addr[59345]= 1000068799;
assign addr[59346]= 931758235;
assign addr[59347]= 862265664;
assign addr[59348]= 791679244;
assign addr[59349]= 720088517;
assign addr[59350]= 647584304;
assign addr[59351]= 574258580;
assign addr[59352]= 500204365;
assign addr[59353]= 425515602;
assign addr[59354]= 350287041;
assign addr[59355]= 274614114;
assign addr[59356]= 198592817;
assign addr[59357]= 122319591;
assign addr[59358]= 45891193;
assign addr[59359]= -30595422;
assign addr[59360]= -107043224;
assign addr[59361]= -183355234;
assign addr[59362]= -259434643;
assign addr[59363]= -335184940;
assign addr[59364]= -410510029;
assign addr[59365]= -485314355;
assign addr[59366]= -559503022;
assign addr[59367]= -632981917;
assign addr[59368]= -705657826;
assign addr[59369]= -777438554;
assign addr[59370]= -848233042;
assign addr[59371]= -917951481;
assign addr[59372]= -986505429;
assign addr[59373]= -1053807919;
assign addr[59374]= -1119773573;
assign addr[59375]= -1184318708;
assign addr[59376]= -1247361445;
assign addr[59377]= -1308821808;
assign addr[59378]= -1368621831;
assign addr[59379]= -1426685652;
assign addr[59380]= -1482939614;
assign addr[59381]= -1537312353;
assign addr[59382]= -1589734894;
assign addr[59383]= -1640140734;
assign addr[59384]= -1688465931;
assign addr[59385]= -1734649179;
assign addr[59386]= -1778631892;
assign addr[59387]= -1820358275;
assign addr[59388]= -1859775393;
assign addr[59389]= -1896833245;
assign addr[59390]= -1931484818;
assign addr[59391]= -1963686155;
assign addr[59392]= -1993396407;
assign addr[59393]= -2020577882;
assign addr[59394]= -2045196100;
assign addr[59395]= -2067219829;
assign addr[59396]= -2086621133;
assign addr[59397]= -2103375398;
assign addr[59398]= -2117461370;
assign addr[59399]= -2128861181;
assign addr[59400]= -2137560369;
assign addr[59401]= -2143547897;
assign addr[59402]= -2146816171;
assign addr[59403]= -2147361045;
assign addr[59404]= -2145181827;
assign addr[59405]= -2140281282;
assign addr[59406]= -2132665626;
assign addr[59407]= -2122344521;
assign addr[59408]= -2109331059;
assign addr[59409]= -2093641749;
assign addr[59410]= -2075296495;
assign addr[59411]= -2054318569;
assign addr[59412]= -2030734582;
assign addr[59413]= -2004574453;
assign addr[59414]= -1975871368;
assign addr[59415]= -1944661739;
assign addr[59416]= -1910985158;
assign addr[59417]= -1874884346;
assign addr[59418]= -1836405100;
assign addr[59419]= -1795596234;
assign addr[59420]= -1752509516;
assign addr[59421]= -1707199606;
assign addr[59422]= -1659723983;
assign addr[59423]= -1610142873;
assign addr[59424]= -1558519173;
assign addr[59425]= -1504918373;
assign addr[59426]= -1449408469;
assign addr[59427]= -1392059879;
assign addr[59428]= -1332945355;
assign addr[59429]= -1272139887;
assign addr[59430]= -1209720613;
assign addr[59431]= -1145766716;
assign addr[59432]= -1080359326;
assign addr[59433]= -1013581418;
assign addr[59434]= -945517704;
assign addr[59435]= -876254528;
assign addr[59436]= -805879757;
assign addr[59437]= -734482665;
assign addr[59438]= -662153826;
assign addr[59439]= -588984994;
assign addr[59440]= -515068990;
assign addr[59441]= -440499581;
assign addr[59442]= -365371365;
assign addr[59443]= -289779648;
assign addr[59444]= -213820322;
assign addr[59445]= -137589750;
assign addr[59446]= -61184634;
assign addr[59447]= 15298099;
assign addr[59448]= 91761426;
assign addr[59449]= 168108346;
assign addr[59450]= 244242007;
assign addr[59451]= 320065829;
assign addr[59452]= 395483624;
assign addr[59453]= 470399716;
assign addr[59454]= 544719071;
assign addr[59455]= 618347408;
assign addr[59456]= 691191324;
assign addr[59457]= 763158411;
assign addr[59458]= 834157373;
assign addr[59459]= 904098143;
assign addr[59460]= 972891995;
assign addr[59461]= 1040451659;
assign addr[59462]= 1106691431;
assign addr[59463]= 1171527280;
assign addr[59464]= 1234876957;
assign addr[59465]= 1296660098;
assign addr[59466]= 1356798326;
assign addr[59467]= 1415215352;
assign addr[59468]= 1471837070;
assign addr[59469]= 1526591649;
assign addr[59470]= 1579409630;
assign addr[59471]= 1630224009;
assign addr[59472]= 1678970324;
assign addr[59473]= 1725586737;
assign addr[59474]= 1770014111;
assign addr[59475]= 1812196087;
assign addr[59476]= 1852079154;
assign addr[59477]= 1889612716;
assign addr[59478]= 1924749160;
assign addr[59479]= 1957443913;
assign addr[59480]= 1987655498;
assign addr[59481]= 2015345591;
assign addr[59482]= 2040479063;
assign addr[59483]= 2063024031;
assign addr[59484]= 2082951896;
assign addr[59485]= 2100237377;
assign addr[59486]= 2114858546;
assign addr[59487]= 2126796855;
assign addr[59488]= 2136037160;
assign addr[59489]= 2142567738;
assign addr[59490]= 2146380306;
assign addr[59491]= 2147470025;
assign addr[59492]= 2145835515;
assign addr[59493]= 2141478848;
assign addr[59494]= 2134405552;
assign addr[59495]= 2124624598;
assign addr[59496]= 2112148396;
assign addr[59497]= 2096992772;
assign addr[59498]= 2079176953;
assign addr[59499]= 2058723538;
assign addr[59500]= 2035658475;
assign addr[59501]= 2010011024;
assign addr[59502]= 1981813720;
assign addr[59503]= 1951102334;
assign addr[59504]= 1917915825;
assign addr[59505]= 1882296293;
assign addr[59506]= 1844288924;
assign addr[59507]= 1803941934;
assign addr[59508]= 1761306505;
assign addr[59509]= 1716436725;
assign addr[59510]= 1669389513;
assign addr[59511]= 1620224553;
assign addr[59512]= 1569004214;
assign addr[59513]= 1515793473;
assign addr[59514]= 1460659832;
assign addr[59515]= 1403673233;
assign addr[59516]= 1344905966;
assign addr[59517]= 1284432584;
assign addr[59518]= 1222329801;
assign addr[59519]= 1158676398;
assign addr[59520]= 1093553126;
assign addr[59521]= 1027042599;
assign addr[59522]= 959229189;
assign addr[59523]= 890198924;
assign addr[59524]= 820039373;
assign addr[59525]= 748839539;
assign addr[59526]= 676689746;
assign addr[59527]= 603681519;
assign addr[59528]= 529907477;
assign addr[59529]= 455461206;
assign addr[59530]= 380437148;
assign addr[59531]= 304930476;
assign addr[59532]= 229036977;
assign addr[59533]= 152852926;
assign addr[59534]= 76474970;
assign addr[59535]= 0;
assign addr[59536]= -76474970;
assign addr[59537]= -152852926;
assign addr[59538]= -229036977;
assign addr[59539]= -304930476;
assign addr[59540]= -380437148;
assign addr[59541]= -455461206;
assign addr[59542]= -529907477;
assign addr[59543]= -603681519;
assign addr[59544]= -676689746;
assign addr[59545]= -748839539;
assign addr[59546]= -820039373;
assign addr[59547]= -890198924;
assign addr[59548]= -959229189;
assign addr[59549]= -1027042599;
assign addr[59550]= -1093553126;
assign addr[59551]= -1158676398;
assign addr[59552]= -1222329801;
assign addr[59553]= -1284432584;
assign addr[59554]= -1344905966;
assign addr[59555]= -1403673233;
assign addr[59556]= -1460659832;
assign addr[59557]= -1515793473;
assign addr[59558]= -1569004214;
assign addr[59559]= -1620224553;
assign addr[59560]= -1669389513;
assign addr[59561]= -1716436725;
assign addr[59562]= -1761306505;
assign addr[59563]= -1803941934;
assign addr[59564]= -1844288924;
assign addr[59565]= -1882296293;
assign addr[59566]= -1917915825;
assign addr[59567]= -1951102334;
assign addr[59568]= -1981813720;
assign addr[59569]= -2010011024;
assign addr[59570]= -2035658475;
assign addr[59571]= -2058723538;
assign addr[59572]= -2079176953;
assign addr[59573]= -2096992772;
assign addr[59574]= -2112148396;
assign addr[59575]= -2124624598;
assign addr[59576]= -2134405552;
assign addr[59577]= -2141478848;
assign addr[59578]= -2145835515;
assign addr[59579]= -2147470025;
assign addr[59580]= -2146380306;
assign addr[59581]= -2142567738;
assign addr[59582]= -2136037160;
assign addr[59583]= -2126796855;
assign addr[59584]= -2114858546;
assign addr[59585]= -2100237377;
assign addr[59586]= -2082951896;
assign addr[59587]= -2063024031;
assign addr[59588]= -2040479063;
assign addr[59589]= -2015345591;
assign addr[59590]= -1987655498;
assign addr[59591]= -1957443913;
assign addr[59592]= -1924749160;
assign addr[59593]= -1889612716;
assign addr[59594]= -1852079154;
assign addr[59595]= -1812196087;
assign addr[59596]= -1770014111;
assign addr[59597]= -1725586737;
assign addr[59598]= -1678970324;
assign addr[59599]= -1630224009;
assign addr[59600]= -1579409630;
assign addr[59601]= -1526591649;
assign addr[59602]= -1471837070;
assign addr[59603]= -1415215352;
assign addr[59604]= -1356798326;
assign addr[59605]= -1296660098;
assign addr[59606]= -1234876957;
assign addr[59607]= -1171527280;
assign addr[59608]= -1106691431;
assign addr[59609]= -1040451659;
assign addr[59610]= -972891995;
assign addr[59611]= -904098143;
assign addr[59612]= -834157373;
assign addr[59613]= -763158411;
assign addr[59614]= -691191324;
assign addr[59615]= -618347408;
assign addr[59616]= -544719071;
assign addr[59617]= -470399716;
assign addr[59618]= -395483624;
assign addr[59619]= -320065829;
assign addr[59620]= -244242007;
assign addr[59621]= -168108346;
assign addr[59622]= -91761426;
assign addr[59623]= -15298099;
assign addr[59624]= 61184634;
assign addr[59625]= 137589750;
assign addr[59626]= 213820322;
assign addr[59627]= 289779648;
assign addr[59628]= 365371365;
assign addr[59629]= 440499581;
assign addr[59630]= 515068990;
assign addr[59631]= 588984994;
assign addr[59632]= 662153826;
assign addr[59633]= 734482665;
assign addr[59634]= 805879757;
assign addr[59635]= 876254528;
assign addr[59636]= 945517704;
assign addr[59637]= 1013581418;
assign addr[59638]= 1080359326;
assign addr[59639]= 1145766716;
assign addr[59640]= 1209720613;
assign addr[59641]= 1272139887;
assign addr[59642]= 1332945355;
assign addr[59643]= 1392059879;
assign addr[59644]= 1449408469;
assign addr[59645]= 1504918373;
assign addr[59646]= 1558519173;
assign addr[59647]= 1610142873;
assign addr[59648]= 1659723983;
assign addr[59649]= 1707199606;
assign addr[59650]= 1752509516;
assign addr[59651]= 1795596234;
assign addr[59652]= 1836405100;
assign addr[59653]= 1874884346;
assign addr[59654]= 1910985158;
assign addr[59655]= 1944661739;
assign addr[59656]= 1975871368;
assign addr[59657]= 2004574453;
assign addr[59658]= 2030734582;
assign addr[59659]= 2054318569;
assign addr[59660]= 2075296495;
assign addr[59661]= 2093641749;
assign addr[59662]= 2109331059;
assign addr[59663]= 2122344521;
assign addr[59664]= 2132665626;
assign addr[59665]= 2140281282;
assign addr[59666]= 2145181827;
assign addr[59667]= 2147361045;
assign addr[59668]= 2146816171;
assign addr[59669]= 2143547897;
assign addr[59670]= 2137560369;
assign addr[59671]= 2128861181;
assign addr[59672]= 2117461370;
assign addr[59673]= 2103375398;
assign addr[59674]= 2086621133;
assign addr[59675]= 2067219829;
assign addr[59676]= 2045196100;
assign addr[59677]= 2020577882;
assign addr[59678]= 1993396407;
assign addr[59679]= 1963686155;
assign addr[59680]= 1931484818;
assign addr[59681]= 1896833245;
assign addr[59682]= 1859775393;
assign addr[59683]= 1820358275;
assign addr[59684]= 1778631892;
assign addr[59685]= 1734649179;
assign addr[59686]= 1688465931;
assign addr[59687]= 1640140734;
assign addr[59688]= 1589734894;
assign addr[59689]= 1537312353;
assign addr[59690]= 1482939614;
assign addr[59691]= 1426685652;
assign addr[59692]= 1368621831;
assign addr[59693]= 1308821808;
assign addr[59694]= 1247361445;
assign addr[59695]= 1184318708;
assign addr[59696]= 1119773573;
assign addr[59697]= 1053807919;
assign addr[59698]= 986505429;
assign addr[59699]= 917951481;
assign addr[59700]= 848233042;
assign addr[59701]= 777438554;
assign addr[59702]= 705657826;
assign addr[59703]= 632981917;
assign addr[59704]= 559503022;
assign addr[59705]= 485314355;
assign addr[59706]= 410510029;
assign addr[59707]= 335184940;
assign addr[59708]= 259434643;
assign addr[59709]= 183355234;
assign addr[59710]= 107043224;
assign addr[59711]= 30595422;
assign addr[59712]= -45891193;
assign addr[59713]= -122319591;
assign addr[59714]= -198592817;
assign addr[59715]= -274614114;
assign addr[59716]= -350287041;
assign addr[59717]= -425515602;
assign addr[59718]= -500204365;
assign addr[59719]= -574258580;
assign addr[59720]= -647584304;
assign addr[59721]= -720088517;
assign addr[59722]= -791679244;
assign addr[59723]= -862265664;
assign addr[59724]= -931758235;
assign addr[59725]= -1000068799;
assign addr[59726]= -1067110699;
assign addr[59727]= -1132798888;
assign addr[59728]= -1197050035;
assign addr[59729]= -1259782632;
assign addr[59730]= -1320917099;
assign addr[59731]= -1380375881;
assign addr[59732]= -1438083551;
assign addr[59733]= -1493966902;
assign addr[59734]= -1547955041;
assign addr[59735]= -1599979481;
assign addr[59736]= -1649974225;
assign addr[59737]= -1697875851;
assign addr[59738]= -1743623590;
assign addr[59739]= -1787159411;
assign addr[59740]= -1828428082;
assign addr[59741]= -1867377253;
assign addr[59742]= -1903957513;
assign addr[59743]= -1938122457;
assign addr[59744]= -1969828744;
assign addr[59745]= -1999036154;
assign addr[59746]= -2025707632;
assign addr[59747]= -2049809346;
assign addr[59748]= -2071310720;
assign addr[59749]= -2090184478;
assign addr[59750]= -2106406677;
assign addr[59751]= -2119956737;
assign addr[59752]= -2130817471;
assign addr[59753]= -2138975100;
assign addr[59754]= -2144419275;
assign addr[59755]= -2147143090;
assign addr[59756]= -2147143090;
assign addr[59757]= -2144419275;
assign addr[59758]= -2138975100;
assign addr[59759]= -2130817471;
assign addr[59760]= -2119956737;
assign addr[59761]= -2106406677;
assign addr[59762]= -2090184478;
assign addr[59763]= -2071310720;
assign addr[59764]= -2049809346;
assign addr[59765]= -2025707632;
assign addr[59766]= -1999036154;
assign addr[59767]= -1969828744;
assign addr[59768]= -1938122457;
assign addr[59769]= -1903957513;
assign addr[59770]= -1867377253;
assign addr[59771]= -1828428082;
assign addr[59772]= -1787159411;
assign addr[59773]= -1743623590;
assign addr[59774]= -1697875851;
assign addr[59775]= -1649974225;
assign addr[59776]= -1599979481;
assign addr[59777]= -1547955041;
assign addr[59778]= -1493966902;
assign addr[59779]= -1438083551;
assign addr[59780]= -1380375881;
assign addr[59781]= -1320917099;
assign addr[59782]= -1259782632;
assign addr[59783]= -1197050035;
assign addr[59784]= -1132798888;
assign addr[59785]= -1067110699;
assign addr[59786]= -1000068799;
assign addr[59787]= -931758235;
assign addr[59788]= -862265664;
assign addr[59789]= -791679244;
assign addr[59790]= -720088517;
assign addr[59791]= -647584304;
assign addr[59792]= -574258580;
assign addr[59793]= -500204365;
assign addr[59794]= -425515602;
assign addr[59795]= -350287041;
assign addr[59796]= -274614114;
assign addr[59797]= -198592817;
assign addr[59798]= -122319591;
assign addr[59799]= -45891193;
assign addr[59800]= 30595422;
assign addr[59801]= 107043224;
assign addr[59802]= 183355234;
assign addr[59803]= 259434643;
assign addr[59804]= 335184940;
assign addr[59805]= 410510029;
assign addr[59806]= 485314355;
assign addr[59807]= 559503022;
assign addr[59808]= 632981917;
assign addr[59809]= 705657826;
assign addr[59810]= 777438554;
assign addr[59811]= 848233042;
assign addr[59812]= 917951481;
assign addr[59813]= 986505429;
assign addr[59814]= 1053807919;
assign addr[59815]= 1119773573;
assign addr[59816]= 1184318708;
assign addr[59817]= 1247361445;
assign addr[59818]= 1308821808;
assign addr[59819]= 1368621831;
assign addr[59820]= 1426685652;
assign addr[59821]= 1482939614;
assign addr[59822]= 1537312353;
assign addr[59823]= 1589734894;
assign addr[59824]= 1640140734;
assign addr[59825]= 1688465931;
assign addr[59826]= 1734649179;
assign addr[59827]= 1778631892;
assign addr[59828]= 1820358275;
assign addr[59829]= 1859775393;
assign addr[59830]= 1896833245;
assign addr[59831]= 1931484818;
assign addr[59832]= 1963686155;
assign addr[59833]= 1993396407;
assign addr[59834]= 2020577882;
assign addr[59835]= 2045196100;
assign addr[59836]= 2067219829;
assign addr[59837]= 2086621133;
assign addr[59838]= 2103375398;
assign addr[59839]= 2117461370;
assign addr[59840]= 2128861181;
assign addr[59841]= 2137560369;
assign addr[59842]= 2143547897;
assign addr[59843]= 2146816171;
assign addr[59844]= 2147361045;
assign addr[59845]= 2145181827;
assign addr[59846]= 2140281282;
assign addr[59847]= 2132665626;
assign addr[59848]= 2122344521;
assign addr[59849]= 2109331059;
assign addr[59850]= 2093641749;
assign addr[59851]= 2075296495;
assign addr[59852]= 2054318569;
assign addr[59853]= 2030734582;
assign addr[59854]= 2004574453;
assign addr[59855]= 1975871368;
assign addr[59856]= 1944661739;
assign addr[59857]= 1910985158;
assign addr[59858]= 1874884346;
assign addr[59859]= 1836405100;
assign addr[59860]= 1795596234;
assign addr[59861]= 1752509516;
assign addr[59862]= 1707199606;
assign addr[59863]= 1659723983;
assign addr[59864]= 1610142873;
assign addr[59865]= 1558519173;
assign addr[59866]= 1504918373;
assign addr[59867]= 1449408469;
assign addr[59868]= 1392059879;
assign addr[59869]= 1332945355;
assign addr[59870]= 1272139887;
assign addr[59871]= 1209720613;
assign addr[59872]= 1145766716;
assign addr[59873]= 1080359326;
assign addr[59874]= 1013581418;
assign addr[59875]= 945517704;
assign addr[59876]= 876254528;
assign addr[59877]= 805879757;
assign addr[59878]= 734482665;
assign addr[59879]= 662153826;
assign addr[59880]= 588984994;
assign addr[59881]= 515068990;
assign addr[59882]= 440499581;
assign addr[59883]= 365371365;
assign addr[59884]= 289779648;
assign addr[59885]= 213820322;
assign addr[59886]= 137589750;
assign addr[59887]= 61184634;
assign addr[59888]= -15298099;
assign addr[59889]= -91761426;
assign addr[59890]= -168108346;
assign addr[59891]= -244242007;
assign addr[59892]= -320065829;
assign addr[59893]= -395483624;
assign addr[59894]= -470399716;
assign addr[59895]= -544719071;
assign addr[59896]= -618347408;
assign addr[59897]= -691191324;
assign addr[59898]= -763158411;
assign addr[59899]= -834157373;
assign addr[59900]= -904098143;
assign addr[59901]= -972891995;
assign addr[59902]= -1040451659;
assign addr[59903]= -1106691431;
assign addr[59904]= -1171527280;
assign addr[59905]= -1234876957;
assign addr[59906]= -1296660098;
assign addr[59907]= -1356798326;
assign addr[59908]= -1415215352;
assign addr[59909]= -1471837070;
assign addr[59910]= -1526591649;
assign addr[59911]= -1579409630;
assign addr[59912]= -1630224009;
assign addr[59913]= -1678970324;
assign addr[59914]= -1725586737;
assign addr[59915]= -1770014111;
assign addr[59916]= -1812196087;
assign addr[59917]= -1852079154;
assign addr[59918]= -1889612716;
assign addr[59919]= -1924749160;
assign addr[59920]= -1957443913;
assign addr[59921]= -1987655498;
assign addr[59922]= -2015345591;
assign addr[59923]= -2040479063;
assign addr[59924]= -2063024031;
assign addr[59925]= -2082951896;
assign addr[59926]= -2100237377;
assign addr[59927]= -2114858546;
assign addr[59928]= -2126796855;
assign addr[59929]= -2136037160;
assign addr[59930]= -2142567738;
assign addr[59931]= -2146380306;
assign addr[59932]= -2147470025;
assign addr[59933]= -2145835515;
assign addr[59934]= -2141478848;
assign addr[59935]= -2134405552;
assign addr[59936]= -2124624598;
assign addr[59937]= -2112148396;
assign addr[59938]= -2096992772;
assign addr[59939]= -2079176953;
assign addr[59940]= -2058723538;
assign addr[59941]= -2035658475;
assign addr[59942]= -2010011024;
assign addr[59943]= -1981813720;
assign addr[59944]= -1951102334;
assign addr[59945]= -1917915825;
assign addr[59946]= -1882296293;
assign addr[59947]= -1844288924;
assign addr[59948]= -1803941934;
assign addr[59949]= -1761306505;
assign addr[59950]= -1716436725;
assign addr[59951]= -1669389513;
assign addr[59952]= -1620224553;
assign addr[59953]= -1569004214;
assign addr[59954]= -1515793473;
assign addr[59955]= -1460659832;
assign addr[59956]= -1403673233;
assign addr[59957]= -1344905966;
assign addr[59958]= -1284432584;
assign addr[59959]= -1222329801;
assign addr[59960]= -1158676398;
assign addr[59961]= -1093553126;
assign addr[59962]= -1027042599;
assign addr[59963]= -959229189;
assign addr[59964]= -890198924;
assign addr[59965]= -820039373;
assign addr[59966]= -748839539;
assign addr[59967]= -676689746;
assign addr[59968]= -603681519;
assign addr[59969]= -529907477;
assign addr[59970]= -455461206;
assign addr[59971]= -380437148;
assign addr[59972]= -304930476;
assign addr[59973]= -229036977;
assign addr[59974]= -152852926;
assign addr[59975]= -76474970;
assign addr[59976]= 0;
assign addr[59977]= 76474970;
assign addr[59978]= 152852926;
assign addr[59979]= 229036977;
assign addr[59980]= 304930476;
assign addr[59981]= 380437148;
assign addr[59982]= 455461206;
assign addr[59983]= 529907477;
assign addr[59984]= 603681519;
assign addr[59985]= 676689746;
assign addr[59986]= 748839539;
assign addr[59987]= 820039373;
assign addr[59988]= 890198924;
assign addr[59989]= 959229189;
assign addr[59990]= 1027042599;
assign addr[59991]= 1093553126;
assign addr[59992]= 1158676398;
assign addr[59993]= 1222329801;
assign addr[59994]= 1284432584;
assign addr[59995]= 1344905966;
assign addr[59996]= 1403673233;
assign addr[59997]= 1460659832;
assign addr[59998]= 1515793473;
assign addr[59999]= 1569004214;
assign addr[60000]= 1620224553;
assign addr[60001]= 1669389513;
assign addr[60002]= 1716436725;
assign addr[60003]= 1761306505;
assign addr[60004]= 1803941934;
assign addr[60005]= 1844288924;
assign addr[60006]= 1882296293;
assign addr[60007]= 1917915825;
assign addr[60008]= 1951102334;
assign addr[60009]= 1981813720;
assign addr[60010]= 2010011024;
assign addr[60011]= 2035658475;
assign addr[60012]= 2058723538;
assign addr[60013]= 2079176953;
assign addr[60014]= 2096992772;
assign addr[60015]= 2112148396;
assign addr[60016]= 2124624598;
assign addr[60017]= 2134405552;
assign addr[60018]= 2141478848;
assign addr[60019]= 2145835515;
assign addr[60020]= 2147470025;
assign addr[60021]= 2146380306;
assign addr[60022]= 2142567738;
assign addr[60023]= 2136037160;
assign addr[60024]= 2126796855;
assign addr[60025]= 2114858546;
assign addr[60026]= 2100237377;
assign addr[60027]= 2082951896;
assign addr[60028]= 2063024031;
assign addr[60029]= 2040479063;
assign addr[60030]= 2015345591;
assign addr[60031]= 1987655498;
assign addr[60032]= 1957443913;
assign addr[60033]= 1924749160;
assign addr[60034]= 1889612716;
assign addr[60035]= 1852079154;
assign addr[60036]= 1812196087;
assign addr[60037]= 1770014111;
assign addr[60038]= 1725586737;
assign addr[60039]= 1678970324;
assign addr[60040]= 1630224009;
assign addr[60041]= 1579409630;
assign addr[60042]= 1526591649;
assign addr[60043]= 1471837070;
assign addr[60044]= 1415215352;
assign addr[60045]= 1356798326;
assign addr[60046]= 1296660098;
assign addr[60047]= 1234876957;
assign addr[60048]= 1171527280;
assign addr[60049]= 1106691431;
assign addr[60050]= 1040451659;
assign addr[60051]= 972891995;
assign addr[60052]= 904098143;
assign addr[60053]= 834157373;
assign addr[60054]= 763158411;
assign addr[60055]= 691191324;
assign addr[60056]= 618347408;
assign addr[60057]= 544719071;
assign addr[60058]= 470399716;
assign addr[60059]= 395483624;
assign addr[60060]= 320065829;
assign addr[60061]= 244242007;
assign addr[60062]= 168108346;
assign addr[60063]= 91761426;
assign addr[60064]= 15298099;
assign addr[60065]= -61184634;
assign addr[60066]= -137589750;
assign addr[60067]= -213820322;
assign addr[60068]= -289779648;
assign addr[60069]= -365371365;
assign addr[60070]= -440499581;
assign addr[60071]= -515068990;
assign addr[60072]= -588984994;
assign addr[60073]= -662153826;
assign addr[60074]= -734482665;
assign addr[60075]= -805879757;
assign addr[60076]= -876254528;
assign addr[60077]= -945517704;
assign addr[60078]= -1013581418;
assign addr[60079]= -1080359326;
assign addr[60080]= -1145766716;
assign addr[60081]= -1209720613;
assign addr[60082]= -1272139887;
assign addr[60083]= -1332945355;
assign addr[60084]= -1392059879;
assign addr[60085]= -1449408469;
assign addr[60086]= -1504918373;
assign addr[60087]= -1558519173;
assign addr[60088]= -1610142873;
assign addr[60089]= -1659723983;
assign addr[60090]= -1707199606;
assign addr[60091]= -1752509516;
assign addr[60092]= -1795596234;
assign addr[60093]= -1836405100;
assign addr[60094]= -1874884346;
assign addr[60095]= -1910985158;
assign addr[60096]= -1944661739;
assign addr[60097]= -1975871368;
assign addr[60098]= -2004574453;
assign addr[60099]= -2030734582;
assign addr[60100]= -2054318569;
assign addr[60101]= -2075296495;
assign addr[60102]= -2093641749;
assign addr[60103]= -2109331059;
assign addr[60104]= -2122344521;
assign addr[60105]= -2132665626;
assign addr[60106]= -2140281282;
assign addr[60107]= -2145181827;
assign addr[60108]= -2147361045;
assign addr[60109]= -2146816171;
assign addr[60110]= -2143547897;
assign addr[60111]= -2137560369;
assign addr[60112]= -2128861181;
assign addr[60113]= -2117461370;
assign addr[60114]= -2103375398;
assign addr[60115]= -2086621133;
assign addr[60116]= -2067219829;
assign addr[60117]= -2045196100;
assign addr[60118]= -2020577882;
assign addr[60119]= -1993396407;
assign addr[60120]= -1963686155;
assign addr[60121]= -1931484818;
assign addr[60122]= -1896833245;
assign addr[60123]= -1859775393;
assign addr[60124]= -1820358275;
assign addr[60125]= -1778631892;
assign addr[60126]= -1734649179;
assign addr[60127]= -1688465931;
assign addr[60128]= -1640140734;
assign addr[60129]= -1589734894;
assign addr[60130]= -1537312353;
assign addr[60131]= -1482939614;
assign addr[60132]= -1426685652;
assign addr[60133]= -1368621831;
assign addr[60134]= -1308821808;
assign addr[60135]= -1247361445;
assign addr[60136]= -1184318708;
assign addr[60137]= -1119773573;
assign addr[60138]= -1053807919;
assign addr[60139]= -986505429;
assign addr[60140]= -917951481;
assign addr[60141]= -848233042;
assign addr[60142]= -777438554;
assign addr[60143]= -705657826;
assign addr[60144]= -632981917;
assign addr[60145]= -559503022;
assign addr[60146]= -485314355;
assign addr[60147]= -410510029;
assign addr[60148]= -335184940;
assign addr[60149]= -259434643;
assign addr[60150]= -183355234;
assign addr[60151]= -107043224;
assign addr[60152]= -30595422;
assign addr[60153]= 45891193;
assign addr[60154]= 122319591;
assign addr[60155]= 198592817;
assign addr[60156]= 274614114;
assign addr[60157]= 350287041;
assign addr[60158]= 425515602;
assign addr[60159]= 500204365;
assign addr[60160]= 574258580;
assign addr[60161]= 647584304;
assign addr[60162]= 720088517;
assign addr[60163]= 791679244;
assign addr[60164]= 862265664;
assign addr[60165]= 931758235;
assign addr[60166]= 1000068799;
assign addr[60167]= 1067110699;
assign addr[60168]= 1132798888;
assign addr[60169]= 1197050035;
assign addr[60170]= 1259782632;
assign addr[60171]= 1320917099;
assign addr[60172]= 1380375881;
assign addr[60173]= 1438083551;
assign addr[60174]= 1493966902;
assign addr[60175]= 1547955041;
assign addr[60176]= 1599979481;
assign addr[60177]= 1649974225;
assign addr[60178]= 1697875851;
assign addr[60179]= 1743623590;
assign addr[60180]= 1787159411;
assign addr[60181]= 1828428082;
assign addr[60182]= 1867377253;
assign addr[60183]= 1903957513;
assign addr[60184]= 1938122457;
assign addr[60185]= 1969828744;
assign addr[60186]= 1999036154;
assign addr[60187]= 2025707632;
assign addr[60188]= 2049809346;
assign addr[60189]= 2071310720;
assign addr[60190]= 2090184478;
assign addr[60191]= 2106406677;
assign addr[60192]= 2119956737;
assign addr[60193]= 2130817471;
assign addr[60194]= 2138975100;
assign addr[60195]= 2144419275;
assign addr[60196]= 2147143090;
assign addr[60197]= 2147143090;
assign addr[60198]= 2144419275;
assign addr[60199]= 2138975100;
assign addr[60200]= 2130817471;
assign addr[60201]= 2119956737;
assign addr[60202]= 2106406677;
assign addr[60203]= 2090184478;
assign addr[60204]= 2071310720;
assign addr[60205]= 2049809346;
assign addr[60206]= 2025707632;
assign addr[60207]= 1999036154;
assign addr[60208]= 1969828744;
assign addr[60209]= 1938122457;
assign addr[60210]= 1903957513;
assign addr[60211]= 1867377253;
assign addr[60212]= 1828428082;
assign addr[60213]= 1787159411;
assign addr[60214]= 1743623590;
assign addr[60215]= 1697875851;
assign addr[60216]= 1649974225;
assign addr[60217]= 1599979481;
assign addr[60218]= 1547955041;
assign addr[60219]= 1493966902;
assign addr[60220]= 1438083551;
assign addr[60221]= 1380375881;
assign addr[60222]= 1320917099;
assign addr[60223]= 1259782632;
assign addr[60224]= 1197050035;
assign addr[60225]= 1132798888;
assign addr[60226]= 1067110699;
assign addr[60227]= 1000068799;
assign addr[60228]= 931758235;
assign addr[60229]= 862265664;
assign addr[60230]= 791679244;
assign addr[60231]= 720088517;
assign addr[60232]= 647584304;
assign addr[60233]= 574258580;
assign addr[60234]= 500204365;
assign addr[60235]= 425515602;
assign addr[60236]= 350287041;
assign addr[60237]= 274614114;
assign addr[60238]= 198592817;
assign addr[60239]= 122319591;
assign addr[60240]= 45891193;
assign addr[60241]= -30595422;
assign addr[60242]= -107043224;
assign addr[60243]= -183355234;
assign addr[60244]= -259434643;
assign addr[60245]= -335184940;
assign addr[60246]= -410510029;
assign addr[60247]= -485314355;
assign addr[60248]= -559503022;
assign addr[60249]= -632981917;
assign addr[60250]= -705657826;
assign addr[60251]= -777438554;
assign addr[60252]= -848233042;
assign addr[60253]= -917951481;
assign addr[60254]= -986505429;
assign addr[60255]= -1053807919;
assign addr[60256]= -1119773573;
assign addr[60257]= -1184318708;
assign addr[60258]= -1247361445;
assign addr[60259]= -1308821808;
assign addr[60260]= -1368621831;
assign addr[60261]= -1426685652;
assign addr[60262]= -1482939614;
assign addr[60263]= -1537312353;
assign addr[60264]= -1589734894;
assign addr[60265]= -1640140734;
assign addr[60266]= -1688465931;
assign addr[60267]= -1734649179;
assign addr[60268]= -1778631892;
assign addr[60269]= -1820358275;
assign addr[60270]= -1859775393;
assign addr[60271]= -1896833245;
assign addr[60272]= -1931484818;
assign addr[60273]= -1963686155;
assign addr[60274]= -1993396407;
assign addr[60275]= -2020577882;
assign addr[60276]= -2045196100;
assign addr[60277]= -2067219829;
assign addr[60278]= -2086621133;
assign addr[60279]= -2103375398;
assign addr[60280]= -2117461370;
assign addr[60281]= -2128861181;
assign addr[60282]= -2137560369;
assign addr[60283]= -2143547897;
assign addr[60284]= -2146816171;
assign addr[60285]= -2147361045;
assign addr[60286]= -2145181827;
assign addr[60287]= -2140281282;
assign addr[60288]= -2132665626;
assign addr[60289]= -2122344521;
assign addr[60290]= -2109331059;
assign addr[60291]= -2093641749;
assign addr[60292]= -2075296495;
assign addr[60293]= -2054318569;
assign addr[60294]= -2030734582;
assign addr[60295]= -2004574453;
assign addr[60296]= -1975871368;
assign addr[60297]= -1944661739;
assign addr[60298]= -1910985158;
assign addr[60299]= -1874884346;
assign addr[60300]= -1836405100;
assign addr[60301]= -1795596234;
assign addr[60302]= -1752509516;
assign addr[60303]= -1707199606;
assign addr[60304]= -1659723983;
assign addr[60305]= -1610142873;
assign addr[60306]= -1558519173;
assign addr[60307]= -1504918373;
assign addr[60308]= -1449408469;
assign addr[60309]= -1392059879;
assign addr[60310]= -1332945355;
assign addr[60311]= -1272139887;
assign addr[60312]= -1209720613;
assign addr[60313]= -1145766716;
assign addr[60314]= -1080359326;
assign addr[60315]= -1013581418;
assign addr[60316]= -945517704;
assign addr[60317]= -876254528;
assign addr[60318]= -805879757;
assign addr[60319]= -734482665;
assign addr[60320]= -662153826;
assign addr[60321]= -588984994;
assign addr[60322]= -515068990;
assign addr[60323]= -440499581;
assign addr[60324]= -365371365;
assign addr[60325]= -289779648;
assign addr[60326]= -213820322;
assign addr[60327]= -137589750;
assign addr[60328]= -61184634;
assign addr[60329]= 15298099;
assign addr[60330]= 91761426;
assign addr[60331]= 168108346;
assign addr[60332]= 244242007;
assign addr[60333]= 320065829;
assign addr[60334]= 395483624;
assign addr[60335]= 470399716;
assign addr[60336]= 544719071;
assign addr[60337]= 618347408;
assign addr[60338]= 691191324;
assign addr[60339]= 763158411;
assign addr[60340]= 834157373;
assign addr[60341]= 904098143;
assign addr[60342]= 972891995;
assign addr[60343]= 1040451659;
assign addr[60344]= 1106691431;
assign addr[60345]= 1171527280;
assign addr[60346]= 1234876957;
assign addr[60347]= 1296660098;
assign addr[60348]= 1356798326;
assign addr[60349]= 1415215352;
assign addr[60350]= 1471837070;
assign addr[60351]= 1526591649;
assign addr[60352]= 1579409630;
assign addr[60353]= 1630224009;
assign addr[60354]= 1678970324;
assign addr[60355]= 1725586737;
assign addr[60356]= 1770014111;
assign addr[60357]= 1812196087;
assign addr[60358]= 1852079154;
assign addr[60359]= 1889612716;
assign addr[60360]= 1924749160;
assign addr[60361]= 1957443913;
assign addr[60362]= 1987655498;
assign addr[60363]= 2015345591;
assign addr[60364]= 2040479063;
assign addr[60365]= 2063024031;
assign addr[60366]= 2082951896;
assign addr[60367]= 2100237377;
assign addr[60368]= 2114858546;
assign addr[60369]= 2126796855;
assign addr[60370]= 2136037160;
assign addr[60371]= 2142567738;
assign addr[60372]= 2146380306;
assign addr[60373]= 2147470025;
assign addr[60374]= 2145835515;
assign addr[60375]= 2141478848;
assign addr[60376]= 2134405552;
assign addr[60377]= 2124624598;
assign addr[60378]= 2112148396;
assign addr[60379]= 2096992772;
assign addr[60380]= 2079176953;
assign addr[60381]= 2058723538;
assign addr[60382]= 2035658475;
assign addr[60383]= 2010011024;
assign addr[60384]= 1981813720;
assign addr[60385]= 1951102334;
assign addr[60386]= 1917915825;
assign addr[60387]= 1882296293;
assign addr[60388]= 1844288924;
assign addr[60389]= 1803941934;
assign addr[60390]= 1761306505;
assign addr[60391]= 1716436725;
assign addr[60392]= 1669389513;
assign addr[60393]= 1620224553;
assign addr[60394]= 1569004214;
assign addr[60395]= 1515793473;
assign addr[60396]= 1460659832;
assign addr[60397]= 1403673233;
assign addr[60398]= 1344905966;
assign addr[60399]= 1284432584;
assign addr[60400]= 1222329801;
assign addr[60401]= 1158676398;
assign addr[60402]= 1093553126;
assign addr[60403]= 1027042599;
assign addr[60404]= 959229189;
assign addr[60405]= 890198924;
assign addr[60406]= 820039373;
assign addr[60407]= 748839539;
assign addr[60408]= 676689746;
assign addr[60409]= 603681519;
assign addr[60410]= 529907477;
assign addr[60411]= 455461206;
assign addr[60412]= 380437148;
assign addr[60413]= 304930476;
assign addr[60414]= 229036977;
assign addr[60415]= 152852926;
assign addr[60416]= 76474970;
assign addr[60417]= 0;
assign addr[60418]= -76474970;
assign addr[60419]= -152852926;
assign addr[60420]= -229036977;
assign addr[60421]= -304930476;
assign addr[60422]= -380437148;
assign addr[60423]= -455461206;
assign addr[60424]= -529907477;
assign addr[60425]= -603681519;
assign addr[60426]= -676689746;
assign addr[60427]= -748839539;
assign addr[60428]= -820039373;
assign addr[60429]= -890198924;
assign addr[60430]= -959229189;
assign addr[60431]= -1027042599;
assign addr[60432]= -1093553126;
assign addr[60433]= -1158676398;
assign addr[60434]= -1222329801;
assign addr[60435]= -1284432584;
assign addr[60436]= -1344905966;
assign addr[60437]= -1403673233;
assign addr[60438]= -1460659832;
assign addr[60439]= -1515793473;
assign addr[60440]= -1569004214;
assign addr[60441]= -1620224553;
assign addr[60442]= -1669389513;
assign addr[60443]= -1716436725;
assign addr[60444]= -1761306505;
assign addr[60445]= -1803941934;
assign addr[60446]= -1844288924;
assign addr[60447]= -1882296293;
assign addr[60448]= -1917915825;
assign addr[60449]= -1951102334;
assign addr[60450]= -1981813720;
assign addr[60451]= -2010011024;
assign addr[60452]= -2035658475;
assign addr[60453]= -2058723538;
assign addr[60454]= -2079176953;
assign addr[60455]= -2096992772;
assign addr[60456]= -2112148396;
assign addr[60457]= -2124624598;
assign addr[60458]= -2134405552;
assign addr[60459]= -2141478848;
assign addr[60460]= -2145835515;
assign addr[60461]= -2147470025;
assign addr[60462]= -2146380306;
assign addr[60463]= -2142567738;
assign addr[60464]= -2136037160;
assign addr[60465]= -2126796855;
assign addr[60466]= -2114858546;
assign addr[60467]= -2100237377;
assign addr[60468]= -2082951896;
assign addr[60469]= -2063024031;
assign addr[60470]= -2040479063;
assign addr[60471]= -2015345591;
assign addr[60472]= -1987655498;
assign addr[60473]= -1957443913;
assign addr[60474]= -1924749160;
assign addr[60475]= -1889612716;
assign addr[60476]= -1852079154;
assign addr[60477]= -1812196087;
assign addr[60478]= -1770014111;
assign addr[60479]= -1725586737;
assign addr[60480]= -1678970324;
assign addr[60481]= -1630224009;
assign addr[60482]= -1579409630;
assign addr[60483]= -1526591649;
assign addr[60484]= -1471837070;
assign addr[60485]= -1415215352;
assign addr[60486]= -1356798326;
assign addr[60487]= -1296660098;
assign addr[60488]= -1234876957;
assign addr[60489]= -1171527280;
assign addr[60490]= -1106691431;
assign addr[60491]= -1040451659;
assign addr[60492]= -972891995;
assign addr[60493]= -904098143;
assign addr[60494]= -834157373;
assign addr[60495]= -763158411;
assign addr[60496]= -691191324;
assign addr[60497]= -618347408;
assign addr[60498]= -544719071;
assign addr[60499]= -470399716;
assign addr[60500]= -395483624;
assign addr[60501]= -320065829;
assign addr[60502]= -244242007;
assign addr[60503]= -168108346;
assign addr[60504]= -91761426;
assign addr[60505]= -15298099;
assign addr[60506]= 61184634;
assign addr[60507]= 137589750;
assign addr[60508]= 213820322;
assign addr[60509]= 289779648;
assign addr[60510]= 365371365;
assign addr[60511]= 440499581;
assign addr[60512]= 515068990;
assign addr[60513]= 588984994;
assign addr[60514]= 662153826;
assign addr[60515]= 734482665;
assign addr[60516]= 805879757;
assign addr[60517]= 876254528;
assign addr[60518]= 945517704;
assign addr[60519]= 1013581418;
assign addr[60520]= 1080359326;
assign addr[60521]= 1145766716;
assign addr[60522]= 1209720613;
assign addr[60523]= 1272139887;
assign addr[60524]= 1332945355;
assign addr[60525]= 1392059879;
assign addr[60526]= 1449408469;
assign addr[60527]= 1504918373;
assign addr[60528]= 1558519173;
assign addr[60529]= 1610142873;
assign addr[60530]= 1659723983;
assign addr[60531]= 1707199606;
assign addr[60532]= 1752509516;
assign addr[60533]= 1795596234;
assign addr[60534]= 1836405100;
assign addr[60535]= 1874884346;
assign addr[60536]= 1910985158;
assign addr[60537]= 1944661739;
assign addr[60538]= 1975871368;
assign addr[60539]= 2004574453;
assign addr[60540]= 2030734582;
assign addr[60541]= 2054318569;
assign addr[60542]= 2075296495;
assign addr[60543]= 2093641749;
assign addr[60544]= 2109331059;
assign addr[60545]= 2122344521;
assign addr[60546]= 2132665626;
assign addr[60547]= 2140281282;
assign addr[60548]= 2145181827;
assign addr[60549]= 2147361045;
assign addr[60550]= 2146816171;
assign addr[60551]= 2143547897;
assign addr[60552]= 2137560369;
assign addr[60553]= 2128861181;
assign addr[60554]= 2117461370;
assign addr[60555]= 2103375398;
assign addr[60556]= 2086621133;
assign addr[60557]= 2067219829;
assign addr[60558]= 2045196100;
assign addr[60559]= 2020577882;
assign addr[60560]= 1993396407;
assign addr[60561]= 1963686155;
assign addr[60562]= 1931484818;
assign addr[60563]= 1896833245;
assign addr[60564]= 1859775393;
assign addr[60565]= 1820358275;
assign addr[60566]= 1778631892;
assign addr[60567]= 1734649179;
assign addr[60568]= 1688465931;
assign addr[60569]= 1640140734;
assign addr[60570]= 1589734894;
assign addr[60571]= 1537312353;
assign addr[60572]= 1482939614;
assign addr[60573]= 1426685652;
assign addr[60574]= 1368621831;
assign addr[60575]= 1308821808;
assign addr[60576]= 1247361445;
assign addr[60577]= 1184318708;
assign addr[60578]= 1119773573;
assign addr[60579]= 1053807919;
assign addr[60580]= 986505429;
assign addr[60581]= 917951481;
assign addr[60582]= 848233042;
assign addr[60583]= 777438554;
assign addr[60584]= 705657826;
assign addr[60585]= 632981917;
assign addr[60586]= 559503022;
assign addr[60587]= 485314355;
assign addr[60588]= 410510029;
assign addr[60589]= 335184940;
assign addr[60590]= 259434643;
assign addr[60591]= 183355234;
assign addr[60592]= 107043224;
assign addr[60593]= 30595422;
assign addr[60594]= -45891193;
assign addr[60595]= -122319591;
assign addr[60596]= -198592817;
assign addr[60597]= -274614114;
assign addr[60598]= -350287041;
assign addr[60599]= -425515602;
assign addr[60600]= -500204365;
assign addr[60601]= -574258580;
assign addr[60602]= -647584304;
assign addr[60603]= -720088517;
assign addr[60604]= -791679244;
assign addr[60605]= -862265664;
assign addr[60606]= -931758235;
assign addr[60607]= -1000068799;
assign addr[60608]= -1067110699;
assign addr[60609]= -1132798888;
assign addr[60610]= -1197050035;
assign addr[60611]= -1259782632;
assign addr[60612]= -1320917099;
assign addr[60613]= -1380375881;
assign addr[60614]= -1438083551;
assign addr[60615]= -1493966902;
assign addr[60616]= -1547955041;
assign addr[60617]= -1599979481;
assign addr[60618]= -1649974225;
assign addr[60619]= -1697875851;
assign addr[60620]= -1743623590;
assign addr[60621]= -1787159411;
assign addr[60622]= -1828428082;
assign addr[60623]= -1867377253;
assign addr[60624]= -1903957513;
assign addr[60625]= -1938122457;
assign addr[60626]= -1969828744;
assign addr[60627]= -1999036154;
assign addr[60628]= -2025707632;
assign addr[60629]= -2049809346;
assign addr[60630]= -2071310720;
assign addr[60631]= -2090184478;
assign addr[60632]= -2106406677;
assign addr[60633]= -2119956737;
assign addr[60634]= -2130817471;
assign addr[60635]= -2138975100;
assign addr[60636]= -2144419275;
assign addr[60637]= -2147143090;
assign addr[60638]= -2147143090;
assign addr[60639]= -2144419275;
assign addr[60640]= -2138975100;
assign addr[60641]= -2130817471;
assign addr[60642]= -2119956737;
assign addr[60643]= -2106406677;
assign addr[60644]= -2090184478;
assign addr[60645]= -2071310720;
assign addr[60646]= -2049809346;
assign addr[60647]= -2025707632;
assign addr[60648]= -1999036154;
assign addr[60649]= -1969828744;
assign addr[60650]= -1938122457;
assign addr[60651]= -1903957513;
assign addr[60652]= -1867377253;
assign addr[60653]= -1828428082;
assign addr[60654]= -1787159411;
assign addr[60655]= -1743623590;
assign addr[60656]= -1697875851;
assign addr[60657]= -1649974225;
assign addr[60658]= -1599979481;
assign addr[60659]= -1547955041;
assign addr[60660]= -1493966902;
assign addr[60661]= -1438083551;
assign addr[60662]= -1380375881;
assign addr[60663]= -1320917099;
assign addr[60664]= -1259782632;
assign addr[60665]= -1197050035;
assign addr[60666]= -1132798888;
assign addr[60667]= -1067110699;
assign addr[60668]= -1000068799;
assign addr[60669]= -931758235;
assign addr[60670]= -862265664;
assign addr[60671]= -791679244;
assign addr[60672]= -720088517;
assign addr[60673]= -647584304;
assign addr[60674]= -574258580;
assign addr[60675]= -500204365;
assign addr[60676]= -425515602;
assign addr[60677]= -350287041;
assign addr[60678]= -274614114;
assign addr[60679]= -198592817;
assign addr[60680]= -122319591;
assign addr[60681]= -45891193;
assign addr[60682]= 30595422;
assign addr[60683]= 107043224;
assign addr[60684]= 183355234;
assign addr[60685]= 259434643;
assign addr[60686]= 335184940;
assign addr[60687]= 410510029;
assign addr[60688]= 485314355;
assign addr[60689]= 559503022;
assign addr[60690]= 632981917;
assign addr[60691]= 705657826;
assign addr[60692]= 777438554;
assign addr[60693]= 848233042;
assign addr[60694]= 917951481;
assign addr[60695]= 986505429;
assign addr[60696]= 1053807919;
assign addr[60697]= 1119773573;
assign addr[60698]= 1184318708;
assign addr[60699]= 1247361445;
assign addr[60700]= 1308821808;
assign addr[60701]= 1368621831;
assign addr[60702]= 1426685652;
assign addr[60703]= 1482939614;
assign addr[60704]= 1537312353;
assign addr[60705]= 1589734894;
assign addr[60706]= 1640140734;
assign addr[60707]= 1688465931;
assign addr[60708]= 1734649179;
assign addr[60709]= 1778631892;
assign addr[60710]= 1820358275;
assign addr[60711]= 1859775393;
assign addr[60712]= 1896833245;
assign addr[60713]= 1931484818;
assign addr[60714]= 1963686155;
assign addr[60715]= 1993396407;
assign addr[60716]= 2020577882;
assign addr[60717]= 2045196100;
assign addr[60718]= 2067219829;
assign addr[60719]= 2086621133;
assign addr[60720]= 2103375398;
assign addr[60721]= 2117461370;
assign addr[60722]= 2128861181;
assign addr[60723]= 2137560369;
assign addr[60724]= 2143547897;
assign addr[60725]= 2146816171;
assign addr[60726]= 2147361045;
assign addr[60727]= 2145181827;
assign addr[60728]= 2140281282;
assign addr[60729]= 2132665626;
assign addr[60730]= 2122344521;
assign addr[60731]= 2109331059;
assign addr[60732]= 2093641749;
assign addr[60733]= 2075296495;
assign addr[60734]= 2054318569;
assign addr[60735]= 2030734582;
assign addr[60736]= 2004574453;
assign addr[60737]= 1975871368;
assign addr[60738]= 1944661739;
assign addr[60739]= 1910985158;
assign addr[60740]= 1874884346;
assign addr[60741]= 1836405100;
assign addr[60742]= 1795596234;
assign addr[60743]= 1752509516;
assign addr[60744]= 1707199606;
assign addr[60745]= 1659723983;
assign addr[60746]= 1610142873;
assign addr[60747]= 1558519173;
assign addr[60748]= 1504918373;
assign addr[60749]= 1449408469;
assign addr[60750]= 1392059879;
assign addr[60751]= 1332945355;
assign addr[60752]= 1272139887;
assign addr[60753]= 1209720613;
assign addr[60754]= 1145766716;
assign addr[60755]= 1080359326;
assign addr[60756]= 1013581418;
assign addr[60757]= 945517704;
assign addr[60758]= 876254528;
assign addr[60759]= 805879757;
assign addr[60760]= 734482665;
assign addr[60761]= 662153826;
assign addr[60762]= 588984994;
assign addr[60763]= 515068990;
assign addr[60764]= 440499581;
assign addr[60765]= 365371365;
assign addr[60766]= 289779648;
assign addr[60767]= 213820322;
assign addr[60768]= 137589750;
assign addr[60769]= 61184634;
assign addr[60770]= -15298099;
assign addr[60771]= -91761426;
assign addr[60772]= -168108346;
assign addr[60773]= -244242007;
assign addr[60774]= -320065829;
assign addr[60775]= -395483624;
assign addr[60776]= -470399716;
assign addr[60777]= -544719071;
assign addr[60778]= -618347408;
assign addr[60779]= -691191324;
assign addr[60780]= -763158411;
assign addr[60781]= -834157373;
assign addr[60782]= -904098143;
assign addr[60783]= -972891995;
assign addr[60784]= -1040451659;
assign addr[60785]= -1106691431;
assign addr[60786]= -1171527280;
assign addr[60787]= -1234876957;
assign addr[60788]= -1296660098;
assign addr[60789]= -1356798326;
assign addr[60790]= -1415215352;
assign addr[60791]= -1471837070;
assign addr[60792]= -1526591649;
assign addr[60793]= -1579409630;
assign addr[60794]= -1630224009;
assign addr[60795]= -1678970324;
assign addr[60796]= -1725586737;
assign addr[60797]= -1770014111;
assign addr[60798]= -1812196087;
assign addr[60799]= -1852079154;
assign addr[60800]= -1889612716;
assign addr[60801]= -1924749160;
assign addr[60802]= -1957443913;
assign addr[60803]= -1987655498;
assign addr[60804]= -2015345591;
assign addr[60805]= -2040479063;
assign addr[60806]= -2063024031;
assign addr[60807]= -2082951896;
assign addr[60808]= -2100237377;
assign addr[60809]= -2114858546;
assign addr[60810]= -2126796855;
assign addr[60811]= -2136037160;
assign addr[60812]= -2142567738;
assign addr[60813]= -2146380306;
assign addr[60814]= -2147470025;
assign addr[60815]= -2145835515;
assign addr[60816]= -2141478848;
assign addr[60817]= -2134405552;
assign addr[60818]= -2124624598;
assign addr[60819]= -2112148396;
assign addr[60820]= -2096992772;
assign addr[60821]= -2079176953;
assign addr[60822]= -2058723538;
assign addr[60823]= -2035658475;
assign addr[60824]= -2010011024;
assign addr[60825]= -1981813720;
assign addr[60826]= -1951102334;
assign addr[60827]= -1917915825;
assign addr[60828]= -1882296293;
assign addr[60829]= -1844288924;
assign addr[60830]= -1803941934;
assign addr[60831]= -1761306505;
assign addr[60832]= -1716436725;
assign addr[60833]= -1669389513;
assign addr[60834]= -1620224553;
assign addr[60835]= -1569004214;
assign addr[60836]= -1515793473;
assign addr[60837]= -1460659832;
assign addr[60838]= -1403673233;
assign addr[60839]= -1344905966;
assign addr[60840]= -1284432584;
assign addr[60841]= -1222329801;
assign addr[60842]= -1158676398;
assign addr[60843]= -1093553126;
assign addr[60844]= -1027042599;
assign addr[60845]= -959229189;
assign addr[60846]= -890198924;
assign addr[60847]= -820039373;
assign addr[60848]= -748839539;
assign addr[60849]= -676689746;
assign addr[60850]= -603681519;
assign addr[60851]= -529907477;
assign addr[60852]= -455461206;
assign addr[60853]= -380437148;
assign addr[60854]= -304930476;
assign addr[60855]= -229036977;
assign addr[60856]= -152852926;
assign addr[60857]= -76474970;
assign addr[60858]= 0;
assign addr[60859]= 76474970;
assign addr[60860]= 152852926;
assign addr[60861]= 229036977;
assign addr[60862]= 304930476;
assign addr[60863]= 380437148;
assign addr[60864]= 455461206;
assign addr[60865]= 529907477;
assign addr[60866]= 603681519;
assign addr[60867]= 676689746;
assign addr[60868]= 748839539;
assign addr[60869]= 820039373;
assign addr[60870]= 890198924;
assign addr[60871]= 959229189;
assign addr[60872]= 1027042599;
assign addr[60873]= 1093553126;
assign addr[60874]= 1158676398;
assign addr[60875]= 1222329801;
assign addr[60876]= 1284432584;
assign addr[60877]= 1344905966;
assign addr[60878]= 1403673233;
assign addr[60879]= 1460659832;
assign addr[60880]= 1515793473;
assign addr[60881]= 1569004214;
assign addr[60882]= 1620224553;
assign addr[60883]= 1669389513;
assign addr[60884]= 1716436725;
assign addr[60885]= 1761306505;
assign addr[60886]= 1803941934;
assign addr[60887]= 1844288924;
assign addr[60888]= 1882296293;
assign addr[60889]= 1917915825;
assign addr[60890]= 1951102334;
assign addr[60891]= 1981813720;
assign addr[60892]= 2010011024;
assign addr[60893]= 2035658475;
assign addr[60894]= 2058723538;
assign addr[60895]= 2079176953;
assign addr[60896]= 2096992772;
assign addr[60897]= 2112148396;
assign addr[60898]= 2124624598;
assign addr[60899]= 2134405552;
assign addr[60900]= 2141478848;
assign addr[60901]= 2145835515;
assign addr[60902]= 2147470025;
assign addr[60903]= 2146380306;
assign addr[60904]= 2142567738;
assign addr[60905]= 2136037160;
assign addr[60906]= 2126796855;
assign addr[60907]= 2114858546;
assign addr[60908]= 2100237377;
assign addr[60909]= 2082951896;
assign addr[60910]= 2063024031;
assign addr[60911]= 2040479063;
assign addr[60912]= 2015345591;
assign addr[60913]= 1987655498;
assign addr[60914]= 1957443913;
assign addr[60915]= 1924749160;
assign addr[60916]= 1889612716;
assign addr[60917]= 1852079154;
assign addr[60918]= 1812196087;
assign addr[60919]= 1770014111;
assign addr[60920]= 1725586737;
assign addr[60921]= 1678970324;
assign addr[60922]= 1630224009;
assign addr[60923]= 1579409630;
assign addr[60924]= 1526591649;
assign addr[60925]= 1471837070;
assign addr[60926]= 1415215352;
assign addr[60927]= 1356798326;
assign addr[60928]= 1296660098;
assign addr[60929]= 1234876957;
assign addr[60930]= 1171527280;
assign addr[60931]= 1106691431;
assign addr[60932]= 1040451659;
assign addr[60933]= 972891995;
assign addr[60934]= 904098143;
assign addr[60935]= 834157373;
assign addr[60936]= 763158411;
assign addr[60937]= 691191324;
assign addr[60938]= 618347408;
assign addr[60939]= 544719071;
assign addr[60940]= 470399716;
assign addr[60941]= 395483624;
assign addr[60942]= 320065829;
assign addr[60943]= 244242007;
assign addr[60944]= 168108346;
assign addr[60945]= 91761426;
assign addr[60946]= 15298099;
assign addr[60947]= -61184634;
assign addr[60948]= -137589750;
assign addr[60949]= -213820322;
assign addr[60950]= -289779648;
assign addr[60951]= -365371365;
assign addr[60952]= -440499581;
assign addr[60953]= -515068990;
assign addr[60954]= -588984994;
assign addr[60955]= -662153826;
assign addr[60956]= -734482665;
assign addr[60957]= -805879757;
assign addr[60958]= -876254528;
assign addr[60959]= -945517704;
assign addr[60960]= -1013581418;
assign addr[60961]= -1080359326;
assign addr[60962]= -1145766716;
assign addr[60963]= -1209720613;
assign addr[60964]= -1272139887;
assign addr[60965]= -1332945355;
assign addr[60966]= -1392059879;
assign addr[60967]= -1449408469;
assign addr[60968]= -1504918373;
assign addr[60969]= -1558519173;
assign addr[60970]= -1610142873;
assign addr[60971]= -1659723983;
assign addr[60972]= -1707199606;
assign addr[60973]= -1752509516;
assign addr[60974]= -1795596234;
assign addr[60975]= -1836405100;
assign addr[60976]= -1874884346;
assign addr[60977]= -1910985158;
assign addr[60978]= -1944661739;
assign addr[60979]= -1975871368;
assign addr[60980]= -2004574453;
assign addr[60981]= -2030734582;
assign addr[60982]= -2054318569;
assign addr[60983]= -2075296495;
assign addr[60984]= -2093641749;
assign addr[60985]= -2109331059;
assign addr[60986]= -2122344521;
assign addr[60987]= -2132665626;
assign addr[60988]= -2140281282;
assign addr[60989]= -2145181827;
assign addr[60990]= -2147361045;
assign addr[60991]= -2146816171;
assign addr[60992]= -2143547897;
assign addr[60993]= -2137560369;
assign addr[60994]= -2128861181;
assign addr[60995]= -2117461370;
assign addr[60996]= -2103375398;
assign addr[60997]= -2086621133;
assign addr[60998]= -2067219829;
assign addr[60999]= -2045196100;
assign addr[61000]= -2020577882;
assign addr[61001]= -1993396407;
assign addr[61002]= -1963686155;
assign addr[61003]= -1931484818;
assign addr[61004]= -1896833245;
assign addr[61005]= -1859775393;
assign addr[61006]= -1820358275;
assign addr[61007]= -1778631892;
assign addr[61008]= -1734649179;
assign addr[61009]= -1688465931;
assign addr[61010]= -1640140734;
assign addr[61011]= -1589734894;
assign addr[61012]= -1537312353;
assign addr[61013]= -1482939614;
assign addr[61014]= -1426685652;
assign addr[61015]= -1368621831;
assign addr[61016]= -1308821808;
assign addr[61017]= -1247361445;
assign addr[61018]= -1184318708;
assign addr[61019]= -1119773573;
assign addr[61020]= -1053807919;
assign addr[61021]= -986505429;
assign addr[61022]= -917951481;
assign addr[61023]= -848233042;
assign addr[61024]= -777438554;
assign addr[61025]= -705657826;
assign addr[61026]= -632981917;
assign addr[61027]= -559503022;
assign addr[61028]= -485314355;
assign addr[61029]= -410510029;
assign addr[61030]= -335184940;
assign addr[61031]= -259434643;
assign addr[61032]= -183355234;
assign addr[61033]= -107043224;
assign addr[61034]= -30595422;
assign addr[61035]= 45891193;
assign addr[61036]= 122319591;
assign addr[61037]= 198592817;
assign addr[61038]= 274614114;
assign addr[61039]= 350287041;
assign addr[61040]= 425515602;
assign addr[61041]= 500204365;
assign addr[61042]= 574258580;
assign addr[61043]= 647584304;
assign addr[61044]= 720088517;
assign addr[61045]= 791679244;
assign addr[61046]= 862265664;
assign addr[61047]= 931758235;
assign addr[61048]= 1000068799;
assign addr[61049]= 1067110699;
assign addr[61050]= 1132798888;
assign addr[61051]= 1197050035;
assign addr[61052]= 1259782632;
assign addr[61053]= 1320917099;
assign addr[61054]= 1380375881;
assign addr[61055]= 1438083551;
assign addr[61056]= 1493966902;
assign addr[61057]= 1547955041;
assign addr[61058]= 1599979481;
assign addr[61059]= 1649974225;
assign addr[61060]= 1697875851;
assign addr[61061]= 1743623590;
assign addr[61062]= 1787159411;
assign addr[61063]= 1828428082;
assign addr[61064]= 1867377253;
assign addr[61065]= 1903957513;
assign addr[61066]= 1938122457;
assign addr[61067]= 1969828744;
assign addr[61068]= 1999036154;
assign addr[61069]= 2025707632;
assign addr[61070]= 2049809346;
assign addr[61071]= 2071310720;
assign addr[61072]= 2090184478;
assign addr[61073]= 2106406677;
assign addr[61074]= 2119956737;
assign addr[61075]= 2130817471;
assign addr[61076]= 2138975100;
assign addr[61077]= 2144419275;
assign addr[61078]= 2147143090;
assign addr[61079]= 2147143090;
assign addr[61080]= 2144419275;
assign addr[61081]= 2138975100;
assign addr[61082]= 2130817471;
assign addr[61083]= 2119956737;
assign addr[61084]= 2106406677;
assign addr[61085]= 2090184478;
assign addr[61086]= 2071310720;
assign addr[61087]= 2049809346;
assign addr[61088]= 2025707632;
assign addr[61089]= 1999036154;
assign addr[61090]= 1969828744;
assign addr[61091]= 1938122457;
assign addr[61092]= 1903957513;
assign addr[61093]= 1867377253;
assign addr[61094]= 1828428082;
assign addr[61095]= 1787159411;
assign addr[61096]= 1743623590;
assign addr[61097]= 1697875851;
assign addr[61098]= 1649974225;
assign addr[61099]= 1599979481;
assign addr[61100]= 1547955041;
assign addr[61101]= 1493966902;
assign addr[61102]= 1438083551;
assign addr[61103]= 1380375881;
assign addr[61104]= 1320917099;
assign addr[61105]= 1259782632;
assign addr[61106]= 1197050035;
assign addr[61107]= 1132798888;
assign addr[61108]= 1067110699;
assign addr[61109]= 1000068799;
assign addr[61110]= 931758235;
assign addr[61111]= 862265664;
assign addr[61112]= 791679244;
assign addr[61113]= 720088517;
assign addr[61114]= 647584304;
assign addr[61115]= 574258580;
assign addr[61116]= 500204365;
assign addr[61117]= 425515602;
assign addr[61118]= 350287041;
assign addr[61119]= 274614114;
assign addr[61120]= 198592817;
assign addr[61121]= 122319591;
assign addr[61122]= 45891193;
assign addr[61123]= -30595422;
assign addr[61124]= -107043224;
assign addr[61125]= -183355234;
assign addr[61126]= -259434643;
assign addr[61127]= -335184940;
assign addr[61128]= -410510029;
assign addr[61129]= -485314355;
assign addr[61130]= -559503022;
assign addr[61131]= -632981917;
assign addr[61132]= -705657826;
assign addr[61133]= -777438554;
assign addr[61134]= -848233042;
assign addr[61135]= -917951481;
assign addr[61136]= -986505429;
assign addr[61137]= -1053807919;
assign addr[61138]= -1119773573;
assign addr[61139]= -1184318708;
assign addr[61140]= -1247361445;
assign addr[61141]= -1308821808;
assign addr[61142]= -1368621831;
assign addr[61143]= -1426685652;
assign addr[61144]= -1482939614;
assign addr[61145]= -1537312353;
assign addr[61146]= -1589734894;
assign addr[61147]= -1640140734;
assign addr[61148]= -1688465931;
assign addr[61149]= -1734649179;
assign addr[61150]= -1778631892;
assign addr[61151]= -1820358275;
assign addr[61152]= -1859775393;
assign addr[61153]= -1896833245;
assign addr[61154]= -1931484818;
assign addr[61155]= -1963686155;
assign addr[61156]= -1993396407;
assign addr[61157]= -2020577882;
assign addr[61158]= -2045196100;
assign addr[61159]= -2067219829;
assign addr[61160]= -2086621133;
assign addr[61161]= -2103375398;
assign addr[61162]= -2117461370;
assign addr[61163]= -2128861181;
assign addr[61164]= -2137560369;
assign addr[61165]= -2143547897;
assign addr[61166]= -2146816171;
assign addr[61167]= -2147361045;
assign addr[61168]= -2145181827;
assign addr[61169]= -2140281282;
assign addr[61170]= -2132665626;
assign addr[61171]= -2122344521;
assign addr[61172]= -2109331059;
assign addr[61173]= -2093641749;
assign addr[61174]= -2075296495;
assign addr[61175]= -2054318569;
assign addr[61176]= -2030734582;
assign addr[61177]= -2004574453;
assign addr[61178]= -1975871368;
assign addr[61179]= -1944661739;
assign addr[61180]= -1910985158;
assign addr[61181]= -1874884346;
assign addr[61182]= -1836405100;
assign addr[61183]= -1795596234;
assign addr[61184]= -1752509516;
assign addr[61185]= -1707199606;
assign addr[61186]= -1659723983;
assign addr[61187]= -1610142873;
assign addr[61188]= -1558519173;
assign addr[61189]= -1504918373;
assign addr[61190]= -1449408469;
assign addr[61191]= -1392059879;
assign addr[61192]= -1332945355;
assign addr[61193]= -1272139887;
assign addr[61194]= -1209720613;
assign addr[61195]= -1145766716;
assign addr[61196]= -1080359326;
assign addr[61197]= -1013581418;
assign addr[61198]= -945517704;
assign addr[61199]= -876254528;
assign addr[61200]= -805879757;
assign addr[61201]= -734482665;
assign addr[61202]= -662153826;
assign addr[61203]= -588984994;
assign addr[61204]= -515068990;
assign addr[61205]= -440499581;
assign addr[61206]= -365371365;
assign addr[61207]= -289779648;
assign addr[61208]= -213820322;
assign addr[61209]= -137589750;
assign addr[61210]= -61184634;
assign addr[61211]= 15298099;
assign addr[61212]= 91761426;
assign addr[61213]= 168108346;
assign addr[61214]= 244242007;
assign addr[61215]= 320065829;
assign addr[61216]= 395483624;
assign addr[61217]= 470399716;
assign addr[61218]= 544719071;
assign addr[61219]= 618347408;
assign addr[61220]= 691191324;
assign addr[61221]= 763158411;
assign addr[61222]= 834157373;
assign addr[61223]= 904098143;
assign addr[61224]= 972891995;
assign addr[61225]= 1040451659;
assign addr[61226]= 1106691431;
assign addr[61227]= 1171527280;
assign addr[61228]= 1234876957;
assign addr[61229]= 1296660098;
assign addr[61230]= 1356798326;
assign addr[61231]= 1415215352;
assign addr[61232]= 1471837070;
assign addr[61233]= 1526591649;
assign addr[61234]= 1579409630;
assign addr[61235]= 1630224009;
assign addr[61236]= 1678970324;
assign addr[61237]= 1725586737;
assign addr[61238]= 1770014111;
assign addr[61239]= 1812196087;
assign addr[61240]= 1852079154;
assign addr[61241]= 1889612716;
assign addr[61242]= 1924749160;
assign addr[61243]= 1957443913;
assign addr[61244]= 1987655498;
assign addr[61245]= 2015345591;
assign addr[61246]= 2040479063;
assign addr[61247]= 2063024031;
assign addr[61248]= 2082951896;
assign addr[61249]= 2100237377;
assign addr[61250]= 2114858546;
assign addr[61251]= 2126796855;
assign addr[61252]= 2136037160;
assign addr[61253]= 2142567738;
assign addr[61254]= 2146380306;
assign addr[61255]= 2147470025;
assign addr[61256]= 2145835515;
assign addr[61257]= 2141478848;
assign addr[61258]= 2134405552;
assign addr[61259]= 2124624598;
assign addr[61260]= 2112148396;
assign addr[61261]= 2096992772;
assign addr[61262]= 2079176953;
assign addr[61263]= 2058723538;
assign addr[61264]= 2035658475;
assign addr[61265]= 2010011024;
assign addr[61266]= 1981813720;
assign addr[61267]= 1951102334;
assign addr[61268]= 1917915825;
assign addr[61269]= 1882296293;
assign addr[61270]= 1844288924;
assign addr[61271]= 1803941934;
assign addr[61272]= 1761306505;
assign addr[61273]= 1716436725;
assign addr[61274]= 1669389513;
assign addr[61275]= 1620224553;
assign addr[61276]= 1569004214;
assign addr[61277]= 1515793473;
assign addr[61278]= 1460659832;
assign addr[61279]= 1403673233;
assign addr[61280]= 1344905966;
assign addr[61281]= 1284432584;
assign addr[61282]= 1222329801;
assign addr[61283]= 1158676398;
assign addr[61284]= 1093553126;
assign addr[61285]= 1027042599;
assign addr[61286]= 959229189;
assign addr[61287]= 890198924;
assign addr[61288]= 820039373;
assign addr[61289]= 748839539;
assign addr[61290]= 676689746;
assign addr[61291]= 603681519;
assign addr[61292]= 529907477;
assign addr[61293]= 455461206;
assign addr[61294]= 380437148;
assign addr[61295]= 304930476;
assign addr[61296]= 229036977;
assign addr[61297]= 152852926;
assign addr[61298]= 76474970;
assign addr[61299]= 0;
assign addr[61300]= -76474970;
assign addr[61301]= -152852926;
assign addr[61302]= -229036977;
assign addr[61303]= -304930476;
assign addr[61304]= -380437148;
assign addr[61305]= -455461206;
assign addr[61306]= -529907477;
assign addr[61307]= -603681519;
assign addr[61308]= -676689746;
assign addr[61309]= -748839539;
assign addr[61310]= -820039373;
assign addr[61311]= -890198924;
assign addr[61312]= -959229189;
assign addr[61313]= -1027042599;
assign addr[61314]= -1093553126;
assign addr[61315]= -1158676398;
assign addr[61316]= -1222329801;
assign addr[61317]= -1284432584;
assign addr[61318]= -1344905966;
assign addr[61319]= -1403673233;
assign addr[61320]= -1460659832;
assign addr[61321]= -1515793473;
assign addr[61322]= -1569004214;
assign addr[61323]= -1620224553;
assign addr[61324]= -1669389513;
assign addr[61325]= -1716436725;
assign addr[61326]= -1761306505;
assign addr[61327]= -1803941934;
assign addr[61328]= -1844288924;
assign addr[61329]= -1882296293;
assign addr[61330]= -1917915825;
assign addr[61331]= -1951102334;
assign addr[61332]= -1981813720;
assign addr[61333]= -2010011024;
assign addr[61334]= -2035658475;
assign addr[61335]= -2058723538;
assign addr[61336]= -2079176953;
assign addr[61337]= -2096992772;
assign addr[61338]= -2112148396;
assign addr[61339]= -2124624598;
assign addr[61340]= -2134405552;
assign addr[61341]= -2141478848;
assign addr[61342]= -2145835515;
assign addr[61343]= -2147470025;
assign addr[61344]= -2146380306;
assign addr[61345]= -2142567738;
assign addr[61346]= -2136037160;
assign addr[61347]= -2126796855;
assign addr[61348]= -2114858546;
assign addr[61349]= -2100237377;
assign addr[61350]= -2082951896;
assign addr[61351]= -2063024031;
assign addr[61352]= -2040479063;
assign addr[61353]= -2015345591;
assign addr[61354]= -1987655498;
assign addr[61355]= -1957443913;
assign addr[61356]= -1924749160;
assign addr[61357]= -1889612716;
assign addr[61358]= -1852079154;
assign addr[61359]= -1812196087;
assign addr[61360]= -1770014111;
assign addr[61361]= -1725586737;
assign addr[61362]= -1678970324;
assign addr[61363]= -1630224009;
assign addr[61364]= -1579409630;
assign addr[61365]= -1526591649;
assign addr[61366]= -1471837070;
assign addr[61367]= -1415215352;
assign addr[61368]= -1356798326;
assign addr[61369]= -1296660098;
assign addr[61370]= -1234876957;
assign addr[61371]= -1171527280;
assign addr[61372]= -1106691431;
assign addr[61373]= -1040451659;
assign addr[61374]= -972891995;
assign addr[61375]= -904098143;
assign addr[61376]= -834157373;
assign addr[61377]= -763158411;
assign addr[61378]= -691191324;
assign addr[61379]= -618347408;
assign addr[61380]= -544719071;
assign addr[61381]= -470399716;
assign addr[61382]= -395483624;
assign addr[61383]= -320065829;
assign addr[61384]= -244242007;
assign addr[61385]= -168108346;
assign addr[61386]= -91761426;
assign addr[61387]= -15298099;
assign addr[61388]= 61184634;
assign addr[61389]= 137589750;
assign addr[61390]= 213820322;
assign addr[61391]= 289779648;
assign addr[61392]= 365371365;
assign addr[61393]= 440499581;
assign addr[61394]= 515068990;
assign addr[61395]= 588984994;
assign addr[61396]= 662153826;
assign addr[61397]= 734482665;
assign addr[61398]= 805879757;
assign addr[61399]= 876254528;
assign addr[61400]= 945517704;
assign addr[61401]= 1013581418;
assign addr[61402]= 1080359326;
assign addr[61403]= 1145766716;
assign addr[61404]= 1209720613;
assign addr[61405]= 1272139887;
assign addr[61406]= 1332945355;
assign addr[61407]= 1392059879;
assign addr[61408]= 1449408469;
assign addr[61409]= 1504918373;
assign addr[61410]= 1558519173;
assign addr[61411]= 1610142873;
assign addr[61412]= 1659723983;
assign addr[61413]= 1707199606;
assign addr[61414]= 1752509516;
assign addr[61415]= 1795596234;
assign addr[61416]= 1836405100;
assign addr[61417]= 1874884346;
assign addr[61418]= 1910985158;
assign addr[61419]= 1944661739;
assign addr[61420]= 1975871368;
assign addr[61421]= 2004574453;
assign addr[61422]= 2030734582;
assign addr[61423]= 2054318569;
assign addr[61424]= 2075296495;
assign addr[61425]= 2093641749;
assign addr[61426]= 2109331059;
assign addr[61427]= 2122344521;
assign addr[61428]= 2132665626;
assign addr[61429]= 2140281282;
assign addr[61430]= 2145181827;
assign addr[61431]= 2147361045;
assign addr[61432]= 2146816171;
assign addr[61433]= 2143547897;
assign addr[61434]= 2137560369;
assign addr[61435]= 2128861181;
assign addr[61436]= 2117461370;
assign addr[61437]= 2103375398;
assign addr[61438]= 2086621133;
assign addr[61439]= 2067219829;
assign addr[61440]= 2045196100;
assign addr[61441]= 2020577882;
assign addr[61442]= 1993396407;
assign addr[61443]= 1963686155;
assign addr[61444]= 1931484818;
assign addr[61445]= 1896833245;
assign addr[61446]= 1859775393;
assign addr[61447]= 1820358275;
assign addr[61448]= 1778631892;
assign addr[61449]= 1734649179;
assign addr[61450]= 1688465931;
assign addr[61451]= 1640140734;
assign addr[61452]= 1589734894;
assign addr[61453]= 1537312353;
assign addr[61454]= 1482939614;
assign addr[61455]= 1426685652;
assign addr[61456]= 1368621831;
assign addr[61457]= 1308821808;
assign addr[61458]= 1247361445;
assign addr[61459]= 1184318708;
assign addr[61460]= 1119773573;
assign addr[61461]= 1053807919;
assign addr[61462]= 986505429;
assign addr[61463]= 917951481;
assign addr[61464]= 848233042;
assign addr[61465]= 777438554;
assign addr[61466]= 705657826;
assign addr[61467]= 632981917;
assign addr[61468]= 559503022;
assign addr[61469]= 485314355;
assign addr[61470]= 410510029;
assign addr[61471]= 335184940;
assign addr[61472]= 259434643;
assign addr[61473]= 183355234;
assign addr[61474]= 107043224;
assign addr[61475]= 30595422;
assign addr[61476]= -45891193;
assign addr[61477]= -122319591;
assign addr[61478]= -198592817;
assign addr[61479]= -274614114;
assign addr[61480]= -350287041;
assign addr[61481]= -425515602;
assign addr[61482]= -500204365;
assign addr[61483]= -574258580;
assign addr[61484]= -647584304;
assign addr[61485]= -720088517;
assign addr[61486]= -791679244;
assign addr[61487]= -862265664;
assign addr[61488]= -931758235;
assign addr[61489]= -1000068799;
assign addr[61490]= -1067110699;
assign addr[61491]= -1132798888;
assign addr[61492]= -1197050035;
assign addr[61493]= -1259782632;
assign addr[61494]= -1320917099;
assign addr[61495]= -1380375881;
assign addr[61496]= -1438083551;
assign addr[61497]= -1493966902;
assign addr[61498]= -1547955041;
assign addr[61499]= -1599979481;
assign addr[61500]= -1649974225;
assign addr[61501]= -1697875851;
assign addr[61502]= -1743623590;
assign addr[61503]= -1787159411;
assign addr[61504]= -1828428082;
assign addr[61505]= -1867377253;
assign addr[61506]= -1903957513;
assign addr[61507]= -1938122457;
assign addr[61508]= -1969828744;
assign addr[61509]= -1999036154;
assign addr[61510]= -2025707632;
assign addr[61511]= -2049809346;
assign addr[61512]= -2071310720;
assign addr[61513]= -2090184478;
assign addr[61514]= -2106406677;
assign addr[61515]= -2119956737;
assign addr[61516]= -2130817471;
assign addr[61517]= -2138975100;
assign addr[61518]= -2144419275;
assign addr[61519]= -2147143090;
assign addr[61520]= -2147143090;
assign addr[61521]= -2144419275;
assign addr[61522]= -2138975100;
assign addr[61523]= -2130817471;
assign addr[61524]= -2119956737;
assign addr[61525]= -2106406677;
assign addr[61526]= -2090184478;
assign addr[61527]= -2071310720;
assign addr[61528]= -2049809346;
assign addr[61529]= -2025707632;
assign addr[61530]= -1999036154;
assign addr[61531]= -1969828744;
assign addr[61532]= -1938122457;
assign addr[61533]= -1903957513;
assign addr[61534]= -1867377253;
assign addr[61535]= -1828428082;
assign addr[61536]= -1787159411;
assign addr[61537]= -1743623590;
assign addr[61538]= -1697875851;
assign addr[61539]= -1649974225;
assign addr[61540]= -1599979481;
assign addr[61541]= -1547955041;
assign addr[61542]= -1493966902;
assign addr[61543]= -1438083551;
assign addr[61544]= -1380375881;
assign addr[61545]= -1320917099;
assign addr[61546]= -1259782632;
assign addr[61547]= -1197050035;
assign addr[61548]= -1132798888;
assign addr[61549]= -1067110699;
assign addr[61550]= -1000068799;
assign addr[61551]= -931758235;
assign addr[61552]= -862265664;
assign addr[61553]= -791679244;
assign addr[61554]= -720088517;
assign addr[61555]= -647584304;
assign addr[61556]= -574258580;
assign addr[61557]= -500204365;
assign addr[61558]= -425515602;
assign addr[61559]= -350287041;
assign addr[61560]= -274614114;
assign addr[61561]= -198592817;
assign addr[61562]= -122319591;
assign addr[61563]= -45891193;
assign addr[61564]= 30595422;
assign addr[61565]= 107043224;
assign addr[61566]= 183355234;
assign addr[61567]= 259434643;
assign addr[61568]= 335184940;
assign addr[61569]= 410510029;
assign addr[61570]= 485314355;
assign addr[61571]= 559503022;
assign addr[61572]= 632981917;
assign addr[61573]= 705657826;
assign addr[61574]= 777438554;
assign addr[61575]= 848233042;
assign addr[61576]= 917951481;
assign addr[61577]= 986505429;
assign addr[61578]= 1053807919;
assign addr[61579]= 1119773573;
assign addr[61580]= 1184318708;
assign addr[61581]= 1247361445;
assign addr[61582]= 1308821808;
assign addr[61583]= 1368621831;
assign addr[61584]= 1426685652;
assign addr[61585]= 1482939614;
assign addr[61586]= 1537312353;
assign addr[61587]= 1589734894;
assign addr[61588]= 1640140734;
assign addr[61589]= 1688465931;
assign addr[61590]= 1734649179;
assign addr[61591]= 1778631892;
assign addr[61592]= 1820358275;
assign addr[61593]= 1859775393;
assign addr[61594]= 1896833245;
assign addr[61595]= 1931484818;
assign addr[61596]= 1963686155;
assign addr[61597]= 1993396407;
assign addr[61598]= 2020577882;
assign addr[61599]= 2045196100;
assign addr[61600]= 2067219829;
assign addr[61601]= 2086621133;
assign addr[61602]= 2103375398;
assign addr[61603]= 2117461370;
assign addr[61604]= 2128861181;
assign addr[61605]= 2137560369;
assign addr[61606]= 2143547897;
assign addr[61607]= 2146816171;
assign addr[61608]= 2147361045;
assign addr[61609]= 2145181827;
assign addr[61610]= 2140281282;
assign addr[61611]= 2132665626;
assign addr[61612]= 2122344521;
assign addr[61613]= 2109331059;
assign addr[61614]= 2093641749;
assign addr[61615]= 2075296495;
assign addr[61616]= 2054318569;
assign addr[61617]= 2030734582;
assign addr[61618]= 2004574453;
assign addr[61619]= 1975871368;
assign addr[61620]= 1944661739;
assign addr[61621]= 1910985158;
assign addr[61622]= 1874884346;
assign addr[61623]= 1836405100;
assign addr[61624]= 1795596234;
assign addr[61625]= 1752509516;
assign addr[61626]= 1707199606;
assign addr[61627]= 1659723983;
assign addr[61628]= 1610142873;
assign addr[61629]= 1558519173;
assign addr[61630]= 1504918373;
assign addr[61631]= 1449408469;
assign addr[61632]= 1392059879;
assign addr[61633]= 1332945355;
assign addr[61634]= 1272139887;
assign addr[61635]= 1209720613;
assign addr[61636]= 1145766716;
assign addr[61637]= 1080359326;
assign addr[61638]= 1013581418;
assign addr[61639]= 945517704;
assign addr[61640]= 876254528;
assign addr[61641]= 805879757;
assign addr[61642]= 734482665;
assign addr[61643]= 662153826;
assign addr[61644]= 588984994;
assign addr[61645]= 515068990;
assign addr[61646]= 440499581;
assign addr[61647]= 365371365;
assign addr[61648]= 289779648;
assign addr[61649]= 213820322;
assign addr[61650]= 137589750;
assign addr[61651]= 61184634;
assign addr[61652]= -15298099;
assign addr[61653]= -91761426;
assign addr[61654]= -168108346;
assign addr[61655]= -244242007;
assign addr[61656]= -320065829;
assign addr[61657]= -395483624;
assign addr[61658]= -470399716;
assign addr[61659]= -544719071;
assign addr[61660]= -618347408;
assign addr[61661]= -691191324;
assign addr[61662]= -763158411;
assign addr[61663]= -834157373;
assign addr[61664]= -904098143;
assign addr[61665]= -972891995;
assign addr[61666]= -1040451659;
assign addr[61667]= -1106691431;
assign addr[61668]= -1171527280;
assign addr[61669]= -1234876957;
assign addr[61670]= -1296660098;
assign addr[61671]= -1356798326;
assign addr[61672]= -1415215352;
assign addr[61673]= -1471837070;
assign addr[61674]= -1526591649;
assign addr[61675]= -1579409630;
assign addr[61676]= -1630224009;
assign addr[61677]= -1678970324;
assign addr[61678]= -1725586737;
assign addr[61679]= -1770014111;
assign addr[61680]= -1812196087;
assign addr[61681]= -1852079154;
assign addr[61682]= -1889612716;
assign addr[61683]= -1924749160;
assign addr[61684]= -1957443913;
assign addr[61685]= -1987655498;
assign addr[61686]= -2015345591;
assign addr[61687]= -2040479063;
assign addr[61688]= -2063024031;
assign addr[61689]= -2082951896;
assign addr[61690]= -2100237377;
assign addr[61691]= -2114858546;
assign addr[61692]= -2126796855;
assign addr[61693]= -2136037160;
assign addr[61694]= -2142567738;
assign addr[61695]= -2146380306;
assign addr[61696]= -2147470025;
assign addr[61697]= -2145835515;
assign addr[61698]= -2141478848;
assign addr[61699]= -2134405552;
assign addr[61700]= -2124624598;
assign addr[61701]= -2112148396;
assign addr[61702]= -2096992772;
assign addr[61703]= -2079176953;
assign addr[61704]= -2058723538;
assign addr[61705]= -2035658475;
assign addr[61706]= -2010011024;
assign addr[61707]= -1981813720;
assign addr[61708]= -1951102334;
assign addr[61709]= -1917915825;
assign addr[61710]= -1882296293;
assign addr[61711]= -1844288924;
assign addr[61712]= -1803941934;
assign addr[61713]= -1761306505;
assign addr[61714]= -1716436725;
assign addr[61715]= -1669389513;
assign addr[61716]= -1620224553;
assign addr[61717]= -1569004214;
assign addr[61718]= -1515793473;
assign addr[61719]= -1460659832;
assign addr[61720]= -1403673233;
assign addr[61721]= -1344905966;
assign addr[61722]= -1284432584;
assign addr[61723]= -1222329801;
assign addr[61724]= -1158676398;
assign addr[61725]= -1093553126;
assign addr[61726]= -1027042599;
assign addr[61727]= -959229189;
assign addr[61728]= -890198924;
assign addr[61729]= -820039373;
assign addr[61730]= -748839539;
assign addr[61731]= -676689746;
assign addr[61732]= -603681519;
assign addr[61733]= -529907477;
assign addr[61734]= -455461206;
assign addr[61735]= -380437148;
assign addr[61736]= -304930476;
assign addr[61737]= -229036977;
assign addr[61738]= -152852926;
assign addr[61739]= -76474970;
assign addr[61740]= 0;
assign addr[61741]= 76474970;
assign addr[61742]= 152852926;
assign addr[61743]= 229036977;
assign addr[61744]= 304930476;
assign addr[61745]= 380437148;
assign addr[61746]= 455461206;
assign addr[61747]= 529907477;
assign addr[61748]= 603681519;
assign addr[61749]= 676689746;
assign addr[61750]= 748839539;
assign addr[61751]= 820039373;
assign addr[61752]= 890198924;
assign addr[61753]= 959229189;
assign addr[61754]= 1027042599;
assign addr[61755]= 1093553126;
assign addr[61756]= 1158676398;
assign addr[61757]= 1222329801;
assign addr[61758]= 1284432584;
assign addr[61759]= 1344905966;
assign addr[61760]= 1403673233;
assign addr[61761]= 1460659832;
assign addr[61762]= 1515793473;
assign addr[61763]= 1569004214;
assign addr[61764]= 1620224553;
assign addr[61765]= 1669389513;
assign addr[61766]= 1716436725;
assign addr[61767]= 1761306505;
assign addr[61768]= 1803941934;
assign addr[61769]= 1844288924;
assign addr[61770]= 1882296293;
assign addr[61771]= 1917915825;
assign addr[61772]= 1951102334;
assign addr[61773]= 1981813720;
assign addr[61774]= 2010011024;
assign addr[61775]= 2035658475;
assign addr[61776]= 2058723538;
assign addr[61777]= 2079176953;
assign addr[61778]= 2096992772;
assign addr[61779]= 2112148396;
assign addr[61780]= 2124624598;
assign addr[61781]= 2134405552;
assign addr[61782]= 2141478848;
assign addr[61783]= 2145835515;
assign addr[61784]= 2147470025;
assign addr[61785]= 2146380306;
assign addr[61786]= 2142567738;
assign addr[61787]= 2136037160;
assign addr[61788]= 2126796855;
assign addr[61789]= 2114858546;
assign addr[61790]= 2100237377;
assign addr[61791]= 2082951896;
assign addr[61792]= 2063024031;
assign addr[61793]= 2040479063;
assign addr[61794]= 2015345591;
assign addr[61795]= 1987655498;
assign addr[61796]= 1957443913;
assign addr[61797]= 1924749160;
assign addr[61798]= 1889612716;
assign addr[61799]= 1852079154;
assign addr[61800]= 1812196087;
assign addr[61801]= 1770014111;
assign addr[61802]= 1725586737;
assign addr[61803]= 1678970324;
assign addr[61804]= 1630224009;
assign addr[61805]= 1579409630;
assign addr[61806]= 1526591649;
assign addr[61807]= 1471837070;
assign addr[61808]= 1415215352;
assign addr[61809]= 1356798326;
assign addr[61810]= 1296660098;
assign addr[61811]= 1234876957;
assign addr[61812]= 1171527280;
assign addr[61813]= 1106691431;
assign addr[61814]= 1040451659;
assign addr[61815]= 972891995;
assign addr[61816]= 904098143;
assign addr[61817]= 834157373;
assign addr[61818]= 763158411;
assign addr[61819]= 691191324;
assign addr[61820]= 618347408;
assign addr[61821]= 544719071;
assign addr[61822]= 470399716;
assign addr[61823]= 395483624;
assign addr[61824]= 320065829;
assign addr[61825]= 244242007;
assign addr[61826]= 168108346;
assign addr[61827]= 91761426;
assign addr[61828]= 15298099;
assign addr[61829]= -61184634;
assign addr[61830]= -137589750;
assign addr[61831]= -213820322;
assign addr[61832]= -289779648;
assign addr[61833]= -365371365;
assign addr[61834]= -440499581;
assign addr[61835]= -515068990;
assign addr[61836]= -588984994;
assign addr[61837]= -662153826;
assign addr[61838]= -734482665;
assign addr[61839]= -805879757;
assign addr[61840]= -876254528;
assign addr[61841]= -945517704;
assign addr[61842]= -1013581418;
assign addr[61843]= -1080359326;
assign addr[61844]= -1145766716;
assign addr[61845]= -1209720613;
assign addr[61846]= -1272139887;
assign addr[61847]= -1332945355;
assign addr[61848]= -1392059879;
assign addr[61849]= -1449408469;
assign addr[61850]= -1504918373;
assign addr[61851]= -1558519173;
assign addr[61852]= -1610142873;
assign addr[61853]= -1659723983;
assign addr[61854]= -1707199606;
assign addr[61855]= -1752509516;
assign addr[61856]= -1795596234;
assign addr[61857]= -1836405100;
assign addr[61858]= -1874884346;
assign addr[61859]= -1910985158;
assign addr[61860]= -1944661739;
assign addr[61861]= -1975871368;
assign addr[61862]= -2004574453;
assign addr[61863]= -2030734582;
assign addr[61864]= -2054318569;
assign addr[61865]= -2075296495;
assign addr[61866]= -2093641749;
assign addr[61867]= -2109331059;
assign addr[61868]= -2122344521;
assign addr[61869]= -2132665626;
assign addr[61870]= -2140281282;
assign addr[61871]= -2145181827;
assign addr[61872]= -2147361045;
assign addr[61873]= -2146816171;
assign addr[61874]= -2143547897;
assign addr[61875]= -2137560369;
assign addr[61876]= -2128861181;
assign addr[61877]= -2117461370;
assign addr[61878]= -2103375398;
assign addr[61879]= -2086621133;
assign addr[61880]= -2067219829;
assign addr[61881]= -2045196100;
assign addr[61882]= -2020577882;
assign addr[61883]= -1993396407;
assign addr[61884]= -1963686155;
assign addr[61885]= -1931484818;
assign addr[61886]= -1896833245;
assign addr[61887]= -1859775393;
assign addr[61888]= -1820358275;
assign addr[61889]= -1778631892;
assign addr[61890]= -1734649179;
assign addr[61891]= -1688465931;
assign addr[61892]= -1640140734;
assign addr[61893]= -1589734894;
assign addr[61894]= -1537312353;
assign addr[61895]= -1482939614;
assign addr[61896]= -1426685652;
assign addr[61897]= -1368621831;
assign addr[61898]= -1308821808;
assign addr[61899]= -1247361445;
assign addr[61900]= -1184318708;
assign addr[61901]= -1119773573;
assign addr[61902]= -1053807919;
assign addr[61903]= -986505429;
assign addr[61904]= -917951481;
assign addr[61905]= -848233042;
assign addr[61906]= -777438554;
assign addr[61907]= -705657826;
assign addr[61908]= -632981917;
assign addr[61909]= -559503022;
assign addr[61910]= -485314355;
assign addr[61911]= -410510029;
assign addr[61912]= -335184940;
assign addr[61913]= -259434643;
assign addr[61914]= -183355234;
assign addr[61915]= -107043224;
assign addr[61916]= -30595422;
assign addr[61917]= 45891193;
assign addr[61918]= 122319591;
assign addr[61919]= 198592817;
assign addr[61920]= 274614114;
assign addr[61921]= 350287041;
assign addr[61922]= 425515602;
assign addr[61923]= 500204365;
assign addr[61924]= 574258580;
assign addr[61925]= 647584304;
assign addr[61926]= 720088517;
assign addr[61927]= 791679244;
assign addr[61928]= 862265664;
assign addr[61929]= 931758235;
assign addr[61930]= 1000068799;
assign addr[61931]= 1067110699;
assign addr[61932]= 1132798888;
assign addr[61933]= 1197050035;
assign addr[61934]= 1259782632;
assign addr[61935]= 1320917099;
assign addr[61936]= 1380375881;
assign addr[61937]= 1438083551;
assign addr[61938]= 1493966902;
assign addr[61939]= 1547955041;
assign addr[61940]= 1599979481;
assign addr[61941]= 1649974225;
assign addr[61942]= 1697875851;
assign addr[61943]= 1743623590;
assign addr[61944]= 1787159411;
assign addr[61945]= 1828428082;
assign addr[61946]= 1867377253;
assign addr[61947]= 1903957513;
assign addr[61948]= 1938122457;
assign addr[61949]= 1969828744;
assign addr[61950]= 1999036154;
assign addr[61951]= 2025707632;
assign addr[61952]= 2049809346;
assign addr[61953]= 2071310720;
assign addr[61954]= 2090184478;
assign addr[61955]= 2106406677;
assign addr[61956]= 2119956737;
assign addr[61957]= 2130817471;
assign addr[61958]= 2138975100;
assign addr[61959]= 2144419275;
assign addr[61960]= 2147143090;
assign addr[61961]= 2147143090;
assign addr[61962]= 2144419275;
assign addr[61963]= 2138975100;
assign addr[61964]= 2130817471;
assign addr[61965]= 2119956737;
assign addr[61966]= 2106406677;
assign addr[61967]= 2090184478;
assign addr[61968]= 2071310720;
assign addr[61969]= 2049809346;
assign addr[61970]= 2025707632;
assign addr[61971]= 1999036154;
assign addr[61972]= 1969828744;
assign addr[61973]= 1938122457;
assign addr[61974]= 1903957513;
assign addr[61975]= 1867377253;
assign addr[61976]= 1828428082;
assign addr[61977]= 1787159411;
assign addr[61978]= 1743623590;
assign addr[61979]= 1697875851;
assign addr[61980]= 1649974225;
assign addr[61981]= 1599979481;
assign addr[61982]= 1547955041;
assign addr[61983]= 1493966902;
assign addr[61984]= 1438083551;
assign addr[61985]= 1380375881;
assign addr[61986]= 1320917099;
assign addr[61987]= 1259782632;
assign addr[61988]= 1197050035;
assign addr[61989]= 1132798888;
assign addr[61990]= 1067110699;
assign addr[61991]= 1000068799;
assign addr[61992]= 931758235;
assign addr[61993]= 862265664;
assign addr[61994]= 791679244;
assign addr[61995]= 720088517;
assign addr[61996]= 647584304;
assign addr[61997]= 574258580;
assign addr[61998]= 500204365;
assign addr[61999]= 425515602;
assign addr[62000]= 350287041;
assign addr[62001]= 274614114;
assign addr[62002]= 198592817;
assign addr[62003]= 122319591;
assign addr[62004]= 45891193;
assign addr[62005]= -30595422;
assign addr[62006]= -107043224;
assign addr[62007]= -183355234;
assign addr[62008]= -259434643;
assign addr[62009]= -335184940;
assign addr[62010]= -410510029;
assign addr[62011]= -485314355;
assign addr[62012]= -559503022;
assign addr[62013]= -632981917;
assign addr[62014]= -705657826;
assign addr[62015]= -777438554;
assign addr[62016]= -848233042;
assign addr[62017]= -917951481;
assign addr[62018]= -986505429;
assign addr[62019]= -1053807919;
assign addr[62020]= -1119773573;
assign addr[62021]= -1184318708;
assign addr[62022]= -1247361445;
assign addr[62023]= -1308821808;
assign addr[62024]= -1368621831;
assign addr[62025]= -1426685652;
assign addr[62026]= -1482939614;
assign addr[62027]= -1537312353;
assign addr[62028]= -1589734894;
assign addr[62029]= -1640140734;
assign addr[62030]= -1688465931;
assign addr[62031]= -1734649179;
assign addr[62032]= -1778631892;
assign addr[62033]= -1820358275;
assign addr[62034]= -1859775393;
assign addr[62035]= -1896833245;
assign addr[62036]= -1931484818;
assign addr[62037]= -1963686155;
assign addr[62038]= -1993396407;
assign addr[62039]= -2020577882;
assign addr[62040]= -2045196100;
assign addr[62041]= -2067219829;
assign addr[62042]= -2086621133;
assign addr[62043]= -2103375398;
assign addr[62044]= -2117461370;
assign addr[62045]= -2128861181;
assign addr[62046]= -2137560369;
assign addr[62047]= -2143547897;
assign addr[62048]= -2146816171;
assign addr[62049]= -2147361045;
assign addr[62050]= -2145181827;
assign addr[62051]= -2140281282;
assign addr[62052]= -2132665626;
assign addr[62053]= -2122344521;
assign addr[62054]= -2109331059;
assign addr[62055]= -2093641749;
assign addr[62056]= -2075296495;
assign addr[62057]= -2054318569;
assign addr[62058]= -2030734582;
assign addr[62059]= -2004574453;
assign addr[62060]= -1975871368;
assign addr[62061]= -1944661739;
assign addr[62062]= -1910985158;
assign addr[62063]= -1874884346;
assign addr[62064]= -1836405100;
assign addr[62065]= -1795596234;
assign addr[62066]= -1752509516;
assign addr[62067]= -1707199606;
assign addr[62068]= -1659723983;
assign addr[62069]= -1610142873;
assign addr[62070]= -1558519173;
assign addr[62071]= -1504918373;
assign addr[62072]= -1449408469;
assign addr[62073]= -1392059879;
assign addr[62074]= -1332945355;
assign addr[62075]= -1272139887;
assign addr[62076]= -1209720613;
assign addr[62077]= -1145766716;
assign addr[62078]= -1080359326;
assign addr[62079]= -1013581418;
assign addr[62080]= -945517704;
assign addr[62081]= -876254528;
assign addr[62082]= -805879757;
assign addr[62083]= -734482665;
assign addr[62084]= -662153826;
assign addr[62085]= -588984994;
assign addr[62086]= -515068990;
assign addr[62087]= -440499581;
assign addr[62088]= -365371365;
assign addr[62089]= -289779648;
assign addr[62090]= -213820322;
assign addr[62091]= -137589750;
assign addr[62092]= -61184634;
assign addr[62093]= 15298099;
assign addr[62094]= 91761426;
assign addr[62095]= 168108346;
assign addr[62096]= 244242007;
assign addr[62097]= 320065829;
assign addr[62098]= 395483624;
assign addr[62099]= 470399716;
assign addr[62100]= 544719071;
assign addr[62101]= 618347408;
assign addr[62102]= 691191324;
assign addr[62103]= 763158411;
assign addr[62104]= 834157373;
assign addr[62105]= 904098143;
assign addr[62106]= 972891995;
assign addr[62107]= 1040451659;
assign addr[62108]= 1106691431;
assign addr[62109]= 1171527280;
assign addr[62110]= 1234876957;
assign addr[62111]= 1296660098;
assign addr[62112]= 1356798326;
assign addr[62113]= 1415215352;
assign addr[62114]= 1471837070;
assign addr[62115]= 1526591649;
assign addr[62116]= 1579409630;
assign addr[62117]= 1630224009;
assign addr[62118]= 1678970324;
assign addr[62119]= 1725586737;
assign addr[62120]= 1770014111;
assign addr[62121]= 1812196087;
assign addr[62122]= 1852079154;
assign addr[62123]= 1889612716;
assign addr[62124]= 1924749160;
assign addr[62125]= 1957443913;
assign addr[62126]= 1987655498;
assign addr[62127]= 2015345591;
assign addr[62128]= 2040479063;
assign addr[62129]= 2063024031;
assign addr[62130]= 2082951896;
assign addr[62131]= 2100237377;
assign addr[62132]= 2114858546;
assign addr[62133]= 2126796855;
assign addr[62134]= 2136037160;
assign addr[62135]= 2142567738;
assign addr[62136]= 2146380306;
assign addr[62137]= 2147470025;
assign addr[62138]= 2145835515;
assign addr[62139]= 2141478848;
assign addr[62140]= 2134405552;
assign addr[62141]= 2124624598;
assign addr[62142]= 2112148396;
assign addr[62143]= 2096992772;
assign addr[62144]= 2079176953;
assign addr[62145]= 2058723538;
assign addr[62146]= 2035658475;
assign addr[62147]= 2010011024;
assign addr[62148]= 1981813720;
assign addr[62149]= 1951102334;
assign addr[62150]= 1917915825;
assign addr[62151]= 1882296293;
assign addr[62152]= 1844288924;
assign addr[62153]= 1803941934;
assign addr[62154]= 1761306505;
assign addr[62155]= 1716436725;
assign addr[62156]= 1669389513;
assign addr[62157]= 1620224553;
assign addr[62158]= 1569004214;
assign addr[62159]= 1515793473;
assign addr[62160]= 1460659832;
assign addr[62161]= 1403673233;
assign addr[62162]= 1344905966;
assign addr[62163]= 1284432584;
assign addr[62164]= 1222329801;
assign addr[62165]= 1158676398;
assign addr[62166]= 1093553126;
assign addr[62167]= 1027042599;
assign addr[62168]= 959229189;
assign addr[62169]= 890198924;
assign addr[62170]= 820039373;
assign addr[62171]= 748839539;
assign addr[62172]= 676689746;
assign addr[62173]= 603681519;
assign addr[62174]= 529907477;
assign addr[62175]= 455461206;
assign addr[62176]= 380437148;
assign addr[62177]= 304930476;
assign addr[62178]= 229036977;
assign addr[62179]= 152852926;
assign addr[62180]= 76474970;
assign addr[62181]= 0;
assign addr[62182]= -76474970;
assign addr[62183]= -152852926;
assign addr[62184]= -229036977;
assign addr[62185]= -304930476;
assign addr[62186]= -380437148;
assign addr[62187]= -455461206;
assign addr[62188]= -529907477;
assign addr[62189]= -603681519;
assign addr[62190]= -676689746;
assign addr[62191]= -748839539;
assign addr[62192]= -820039373;
assign addr[62193]= -890198924;
assign addr[62194]= -959229189;
assign addr[62195]= -1027042599;
assign addr[62196]= -1093553126;
assign addr[62197]= -1158676398;
assign addr[62198]= -1222329801;
assign addr[62199]= -1284432584;
assign addr[62200]= -1344905966;
assign addr[62201]= -1403673233;
assign addr[62202]= -1460659832;
assign addr[62203]= -1515793473;
assign addr[62204]= -1569004214;
assign addr[62205]= -1620224553;
assign addr[62206]= -1669389513;
assign addr[62207]= -1716436725;
assign addr[62208]= -1761306505;
assign addr[62209]= -1803941934;
assign addr[62210]= -1844288924;
assign addr[62211]= -1882296293;
assign addr[62212]= -1917915825;
assign addr[62213]= -1951102334;
assign addr[62214]= -1981813720;
assign addr[62215]= -2010011024;
assign addr[62216]= -2035658475;
assign addr[62217]= -2058723538;
assign addr[62218]= -2079176953;
assign addr[62219]= -2096992772;
assign addr[62220]= -2112148396;
assign addr[62221]= -2124624598;
assign addr[62222]= -2134405552;
assign addr[62223]= -2141478848;
assign addr[62224]= -2145835515;
assign addr[62225]= -2147470025;
assign addr[62226]= -2146380306;
assign addr[62227]= -2142567738;
assign addr[62228]= -2136037160;
assign addr[62229]= -2126796855;
assign addr[62230]= -2114858546;
assign addr[62231]= -2100237377;
assign addr[62232]= -2082951896;
assign addr[62233]= -2063024031;
assign addr[62234]= -2040479063;
assign addr[62235]= -2015345591;
assign addr[62236]= -1987655498;
assign addr[62237]= -1957443913;
assign addr[62238]= -1924749160;
assign addr[62239]= -1889612716;
assign addr[62240]= -1852079154;
assign addr[62241]= -1812196087;
assign addr[62242]= -1770014111;
assign addr[62243]= -1725586737;
assign addr[62244]= -1678970324;
assign addr[62245]= -1630224009;
assign addr[62246]= -1579409630;
assign addr[62247]= -1526591649;
assign addr[62248]= -1471837070;
assign addr[62249]= -1415215352;
assign addr[62250]= -1356798326;
assign addr[62251]= -1296660098;
assign addr[62252]= -1234876957;
assign addr[62253]= -1171527280;
assign addr[62254]= -1106691431;
assign addr[62255]= -1040451659;
assign addr[62256]= -972891995;
assign addr[62257]= -904098143;
assign addr[62258]= -834157373;
assign addr[62259]= -763158411;
assign addr[62260]= -691191324;
assign addr[62261]= -618347408;
assign addr[62262]= -544719071;
assign addr[62263]= -470399716;
assign addr[62264]= -395483624;
assign addr[62265]= -320065829;
assign addr[62266]= -244242007;
assign addr[62267]= -168108346;
assign addr[62268]= -91761426;
assign addr[62269]= -15298099;
assign addr[62270]= 61184634;
assign addr[62271]= 137589750;
assign addr[62272]= 213820322;
assign addr[62273]= 289779648;
assign addr[62274]= 365371365;
assign addr[62275]= 440499581;
assign addr[62276]= 515068990;
assign addr[62277]= 588984994;
assign addr[62278]= 662153826;
assign addr[62279]= 734482665;
assign addr[62280]= 805879757;
assign addr[62281]= 876254528;
assign addr[62282]= 945517704;
assign addr[62283]= 1013581418;
assign addr[62284]= 1080359326;
assign addr[62285]= 1145766716;
assign addr[62286]= 1209720613;
assign addr[62287]= 1272139887;
assign addr[62288]= 1332945355;
assign addr[62289]= 1392059879;
assign addr[62290]= 1449408469;
assign addr[62291]= 1504918373;
assign addr[62292]= 1558519173;
assign addr[62293]= 1610142873;
assign addr[62294]= 1659723983;
assign addr[62295]= 1707199606;
assign addr[62296]= 1752509516;
assign addr[62297]= 1795596234;
assign addr[62298]= 1836405100;
assign addr[62299]= 1874884346;
assign addr[62300]= 1910985158;
assign addr[62301]= 1944661739;
assign addr[62302]= 1975871368;
assign addr[62303]= 2004574453;
assign addr[62304]= 2030734582;
assign addr[62305]= 2054318569;
assign addr[62306]= 2075296495;
assign addr[62307]= 2093641749;
assign addr[62308]= 2109331059;
assign addr[62309]= 2122344521;
assign addr[62310]= 2132665626;
assign addr[62311]= 2140281282;
assign addr[62312]= 2145181827;
assign addr[62313]= 2147361045;
assign addr[62314]= 2146816171;
assign addr[62315]= 2143547897;
assign addr[62316]= 2137560369;
assign addr[62317]= 2128861181;
assign addr[62318]= 2117461370;
assign addr[62319]= 2103375398;
assign addr[62320]= 2086621133;
assign addr[62321]= 2067219829;
assign addr[62322]= 2045196100;
assign addr[62323]= 2020577882;
assign addr[62324]= 1993396407;
assign addr[62325]= 1963686155;
assign addr[62326]= 1931484818;
assign addr[62327]= 1896833245;
assign addr[62328]= 1859775393;
assign addr[62329]= 1820358275;
assign addr[62330]= 1778631892;
assign addr[62331]= 1734649179;
assign addr[62332]= 1688465931;
assign addr[62333]= 1640140734;
assign addr[62334]= 1589734894;
assign addr[62335]= 1537312353;
assign addr[62336]= 1482939614;
assign addr[62337]= 1426685652;
assign addr[62338]= 1368621831;
assign addr[62339]= 1308821808;
assign addr[62340]= 1247361445;
assign addr[62341]= 1184318708;
assign addr[62342]= 1119773573;
assign addr[62343]= 1053807919;
assign addr[62344]= 986505429;
assign addr[62345]= 917951481;
assign addr[62346]= 848233042;
assign addr[62347]= 777438554;
assign addr[62348]= 705657826;
assign addr[62349]= 632981917;
assign addr[62350]= 559503022;
assign addr[62351]= 485314355;
assign addr[62352]= 410510029;
assign addr[62353]= 335184940;
assign addr[62354]= 259434643;
assign addr[62355]= 183355234;
assign addr[62356]= 107043224;
assign addr[62357]= 30595422;
assign addr[62358]= -45891193;
assign addr[62359]= -122319591;
assign addr[62360]= -198592817;
assign addr[62361]= -274614114;
assign addr[62362]= -350287041;
assign addr[62363]= -425515602;
assign addr[62364]= -500204365;
assign addr[62365]= -574258580;
assign addr[62366]= -647584304;
assign addr[62367]= -720088517;
assign addr[62368]= -791679244;
assign addr[62369]= -862265664;
assign addr[62370]= -931758235;
assign addr[62371]= -1000068799;
assign addr[62372]= -1067110699;
assign addr[62373]= -1132798888;
assign addr[62374]= -1197050035;
assign addr[62375]= -1259782632;
assign addr[62376]= -1320917099;
assign addr[62377]= -1380375881;
assign addr[62378]= -1438083551;
assign addr[62379]= -1493966902;
assign addr[62380]= -1547955041;
assign addr[62381]= -1599979481;
assign addr[62382]= -1649974225;
assign addr[62383]= -1697875851;
assign addr[62384]= -1743623590;
assign addr[62385]= -1787159411;
assign addr[62386]= -1828428082;
assign addr[62387]= -1867377253;
assign addr[62388]= -1903957513;
assign addr[62389]= -1938122457;
assign addr[62390]= -1969828744;
assign addr[62391]= -1999036154;
assign addr[62392]= -2025707632;
assign addr[62393]= -2049809346;
assign addr[62394]= -2071310720;
assign addr[62395]= -2090184478;
assign addr[62396]= -2106406677;
assign addr[62397]= -2119956737;
assign addr[62398]= -2130817471;
assign addr[62399]= -2138975100;
assign addr[62400]= -2144419275;
assign addr[62401]= -2147143090;
assign addr[62402]= -2147143090;
assign addr[62403]= -2144419275;
assign addr[62404]= -2138975100;
assign addr[62405]= -2130817471;
assign addr[62406]= -2119956737;
assign addr[62407]= -2106406677;
assign addr[62408]= -2090184478;
assign addr[62409]= -2071310720;
assign addr[62410]= -2049809346;
assign addr[62411]= -2025707632;
assign addr[62412]= -1999036154;
assign addr[62413]= -1969828744;
assign addr[62414]= -1938122457;
assign addr[62415]= -1903957513;
assign addr[62416]= -1867377253;
assign addr[62417]= -1828428082;
assign addr[62418]= -1787159411;
assign addr[62419]= -1743623590;
assign addr[62420]= -1697875851;
assign addr[62421]= -1649974225;
assign addr[62422]= -1599979481;
assign addr[62423]= -1547955041;
assign addr[62424]= -1493966902;
assign addr[62425]= -1438083551;
assign addr[62426]= -1380375881;
assign addr[62427]= -1320917099;
assign addr[62428]= -1259782632;
assign addr[62429]= -1197050035;
assign addr[62430]= -1132798888;
assign addr[62431]= -1067110699;
assign addr[62432]= -1000068799;
assign addr[62433]= -931758235;
assign addr[62434]= -862265664;
assign addr[62435]= -791679244;
assign addr[62436]= -720088517;
assign addr[62437]= -647584304;
assign addr[62438]= -574258580;
assign addr[62439]= -500204365;
assign addr[62440]= -425515602;
assign addr[62441]= -350287041;
assign addr[62442]= -274614114;
assign addr[62443]= -198592817;
assign addr[62444]= -122319591;
assign addr[62445]= -45891193;
assign addr[62446]= 30595422;
assign addr[62447]= 107043224;
assign addr[62448]= 183355234;
assign addr[62449]= 259434643;
assign addr[62450]= 335184940;
assign addr[62451]= 410510029;
assign addr[62452]= 485314355;
assign addr[62453]= 559503022;
assign addr[62454]= 632981917;
assign addr[62455]= 705657826;
assign addr[62456]= 777438554;
assign addr[62457]= 848233042;
assign addr[62458]= 917951481;
assign addr[62459]= 986505429;
assign addr[62460]= 1053807919;
assign addr[62461]= 1119773573;
assign addr[62462]= 1184318708;
assign addr[62463]= 1247361445;
assign addr[62464]= 1308821808;
assign addr[62465]= 1368621831;
assign addr[62466]= 1426685652;
assign addr[62467]= 1482939614;
assign addr[62468]= 1537312353;
assign addr[62469]= 1589734894;
assign addr[62470]= 1640140734;
assign addr[62471]= 1688465931;
assign addr[62472]= 1734649179;
assign addr[62473]= 1778631892;
assign addr[62474]= 1820358275;
assign addr[62475]= 1859775393;
assign addr[62476]= 1896833245;
assign addr[62477]= 1931484818;
assign addr[62478]= 1963686155;
assign addr[62479]= 1993396407;
assign addr[62480]= 2020577882;
assign addr[62481]= 2045196100;
assign addr[62482]= 2067219829;
assign addr[62483]= 2086621133;
assign addr[62484]= 2103375398;
assign addr[62485]= 2117461370;
assign addr[62486]= 2128861181;
assign addr[62487]= 2137560369;
assign addr[62488]= 2143547897;
assign addr[62489]= 2146816171;
assign addr[62490]= 2147361045;
assign addr[62491]= 2145181827;
assign addr[62492]= 2140281282;
assign addr[62493]= 2132665626;
assign addr[62494]= 2122344521;
assign addr[62495]= 2109331059;
assign addr[62496]= 2093641749;
assign addr[62497]= 2075296495;
assign addr[62498]= 2054318569;
assign addr[62499]= 2030734582;
assign addr[62500]= 2004574453;
assign addr[62501]= 1975871368;
assign addr[62502]= 1944661739;
assign addr[62503]= 1910985158;
assign addr[62504]= 1874884346;
assign addr[62505]= 1836405100;
assign addr[62506]= 1795596234;
assign addr[62507]= 1752509516;
assign addr[62508]= 1707199606;
assign addr[62509]= 1659723983;
assign addr[62510]= 1610142873;
assign addr[62511]= 1558519173;
assign addr[62512]= 1504918373;
assign addr[62513]= 1449408469;
assign addr[62514]= 1392059879;
assign addr[62515]= 1332945355;
assign addr[62516]= 1272139887;
assign addr[62517]= 1209720613;
assign addr[62518]= 1145766716;
assign addr[62519]= 1080359326;
assign addr[62520]= 1013581418;
assign addr[62521]= 945517704;
assign addr[62522]= 876254528;
assign addr[62523]= 805879757;
assign addr[62524]= 734482665;
assign addr[62525]= 662153826;
assign addr[62526]= 588984994;
assign addr[62527]= 515068990;
assign addr[62528]= 440499581;
assign addr[62529]= 365371365;
assign addr[62530]= 289779648;
assign addr[62531]= 213820322;
assign addr[62532]= 137589750;
assign addr[62533]= 61184634;
assign addr[62534]= -15298099;
assign addr[62535]= -91761426;
assign addr[62536]= -168108346;
assign addr[62537]= -244242007;
assign addr[62538]= -320065829;
assign addr[62539]= -395483624;
assign addr[62540]= -470399716;
assign addr[62541]= -544719071;
assign addr[62542]= -618347408;
assign addr[62543]= -691191324;
assign addr[62544]= -763158411;
assign addr[62545]= -834157373;
assign addr[62546]= -904098143;
assign addr[62547]= -972891995;
assign addr[62548]= -1040451659;
assign addr[62549]= -1106691431;
assign addr[62550]= -1171527280;
assign addr[62551]= -1234876957;
assign addr[62552]= -1296660098;
assign addr[62553]= -1356798326;
assign addr[62554]= -1415215352;
assign addr[62555]= -1471837070;
assign addr[62556]= -1526591649;
assign addr[62557]= -1579409630;
assign addr[62558]= -1630224009;
assign addr[62559]= -1678970324;
assign addr[62560]= -1725586737;
assign addr[62561]= -1770014111;
assign addr[62562]= -1812196087;
assign addr[62563]= -1852079154;
assign addr[62564]= -1889612716;
assign addr[62565]= -1924749160;
assign addr[62566]= -1957443913;
assign addr[62567]= -1987655498;
assign addr[62568]= -2015345591;
assign addr[62569]= -2040479063;
assign addr[62570]= -2063024031;
assign addr[62571]= -2082951896;
assign addr[62572]= -2100237377;
assign addr[62573]= -2114858546;
assign addr[62574]= -2126796855;
assign addr[62575]= -2136037160;
assign addr[62576]= -2142567738;
assign addr[62577]= -2146380306;
assign addr[62578]= -2147470025;
assign addr[62579]= -2145835515;
assign addr[62580]= -2141478848;
assign addr[62581]= -2134405552;
assign addr[62582]= -2124624598;
assign addr[62583]= -2112148396;
assign addr[62584]= -2096992772;
assign addr[62585]= -2079176953;
assign addr[62586]= -2058723538;
assign addr[62587]= -2035658475;
assign addr[62588]= -2010011024;
assign addr[62589]= -1981813720;
assign addr[62590]= -1951102334;
assign addr[62591]= -1917915825;
assign addr[62592]= -1882296293;
assign addr[62593]= -1844288924;
assign addr[62594]= -1803941934;
assign addr[62595]= -1761306505;
assign addr[62596]= -1716436725;
assign addr[62597]= -1669389513;
assign addr[62598]= -1620224553;
assign addr[62599]= -1569004214;
assign addr[62600]= -1515793473;
assign addr[62601]= -1460659832;
assign addr[62602]= -1403673233;
assign addr[62603]= -1344905966;
assign addr[62604]= -1284432584;
assign addr[62605]= -1222329801;
assign addr[62606]= -1158676398;
assign addr[62607]= -1093553126;
assign addr[62608]= -1027042599;
assign addr[62609]= -959229189;
assign addr[62610]= -890198924;
assign addr[62611]= -820039373;
assign addr[62612]= -748839539;
assign addr[62613]= -676689746;
assign addr[62614]= -603681519;
assign addr[62615]= -529907477;
assign addr[62616]= -455461206;
assign addr[62617]= -380437148;
assign addr[62618]= -304930476;
assign addr[62619]= -229036977;
assign addr[62620]= -152852926;
assign addr[62621]= -76474970;
assign addr[62622]= 0;
assign addr[62623]= 76474970;
assign addr[62624]= 152852926;
assign addr[62625]= 229036977;
assign addr[62626]= 304930476;
assign addr[62627]= 380437148;
assign addr[62628]= 455461206;
assign addr[62629]= 529907477;
assign addr[62630]= 603681519;
assign addr[62631]= 676689746;
assign addr[62632]= 748839539;
assign addr[62633]= 820039373;
assign addr[62634]= 890198924;
assign addr[62635]= 959229189;
assign addr[62636]= 1027042599;
assign addr[62637]= 1093553126;
assign addr[62638]= 1158676398;
assign addr[62639]= 1222329801;
assign addr[62640]= 1284432584;
assign addr[62641]= 1344905966;
assign addr[62642]= 1403673233;
assign addr[62643]= 1460659832;
assign addr[62644]= 1515793473;
assign addr[62645]= 1569004214;
assign addr[62646]= 1620224553;
assign addr[62647]= 1669389513;
assign addr[62648]= 1716436725;
assign addr[62649]= 1761306505;
assign addr[62650]= 1803941934;
assign addr[62651]= 1844288924;
assign addr[62652]= 1882296293;
assign addr[62653]= 1917915825;
assign addr[62654]= 1951102334;
assign addr[62655]= 1981813720;
assign addr[62656]= 2010011024;
assign addr[62657]= 2035658475;
assign addr[62658]= 2058723538;
assign addr[62659]= 2079176953;
assign addr[62660]= 2096992772;
assign addr[62661]= 2112148396;
assign addr[62662]= 2124624598;
assign addr[62663]= 2134405552;
assign addr[62664]= 2141478848;
assign addr[62665]= 2145835515;
assign addr[62666]= 2147470025;
assign addr[62667]= 2146380306;
assign addr[62668]= 2142567738;
assign addr[62669]= 2136037160;
assign addr[62670]= 2126796855;
assign addr[62671]= 2114858546;
assign addr[62672]= 2100237377;
assign addr[62673]= 2082951896;
assign addr[62674]= 2063024031;
assign addr[62675]= 2040479063;
assign addr[62676]= 2015345591;
assign addr[62677]= 1987655498;
assign addr[62678]= 1957443913;
assign addr[62679]= 1924749160;
assign addr[62680]= 1889612716;
assign addr[62681]= 1852079154;
assign addr[62682]= 1812196087;
assign addr[62683]= 1770014111;
assign addr[62684]= 1725586737;
assign addr[62685]= 1678970324;
assign addr[62686]= 1630224009;
assign addr[62687]= 1579409630;
assign addr[62688]= 1526591649;
assign addr[62689]= 1471837070;
assign addr[62690]= 1415215352;
assign addr[62691]= 1356798326;
assign addr[62692]= 1296660098;
assign addr[62693]= 1234876957;
assign addr[62694]= 1171527280;
assign addr[62695]= 1106691431;
assign addr[62696]= 1040451659;
assign addr[62697]= 972891995;
assign addr[62698]= 904098143;
assign addr[62699]= 834157373;
assign addr[62700]= 763158411;
assign addr[62701]= 691191324;
assign addr[62702]= 618347408;
assign addr[62703]= 544719071;
assign addr[62704]= 470399716;
assign addr[62705]= 395483624;
assign addr[62706]= 320065829;
assign addr[62707]= 244242007;
assign addr[62708]= 168108346;
assign addr[62709]= 91761426;
assign addr[62710]= 15298099;
assign addr[62711]= -61184634;
assign addr[62712]= -137589750;
assign addr[62713]= -213820322;
assign addr[62714]= -289779648;
assign addr[62715]= -365371365;
assign addr[62716]= -440499581;
assign addr[62717]= -515068990;
assign addr[62718]= -588984994;
assign addr[62719]= -662153826;
assign addr[62720]= -734482665;
assign addr[62721]= -805879757;
assign addr[62722]= -876254528;
assign addr[62723]= -945517704;
assign addr[62724]= -1013581418;
assign addr[62725]= -1080359326;
assign addr[62726]= -1145766716;
assign addr[62727]= -1209720613;
assign addr[62728]= -1272139887;
assign addr[62729]= -1332945355;
assign addr[62730]= -1392059879;
assign addr[62731]= -1449408469;
assign addr[62732]= -1504918373;
assign addr[62733]= -1558519173;
assign addr[62734]= -1610142873;
assign addr[62735]= -1659723983;
assign addr[62736]= -1707199606;
assign addr[62737]= -1752509516;
assign addr[62738]= -1795596234;
assign addr[62739]= -1836405100;
assign addr[62740]= -1874884346;
assign addr[62741]= -1910985158;
assign addr[62742]= -1944661739;
assign addr[62743]= -1975871368;
assign addr[62744]= -2004574453;
assign addr[62745]= -2030734582;
assign addr[62746]= -2054318569;
assign addr[62747]= -2075296495;
assign addr[62748]= -2093641749;
assign addr[62749]= -2109331059;
assign addr[62750]= -2122344521;
assign addr[62751]= -2132665626;
assign addr[62752]= -2140281282;
assign addr[62753]= -2145181827;
assign addr[62754]= -2147361045;
assign addr[62755]= -2146816171;
assign addr[62756]= -2143547897;
assign addr[62757]= -2137560369;
assign addr[62758]= -2128861181;
assign addr[62759]= -2117461370;
assign addr[62760]= -2103375398;
assign addr[62761]= -2086621133;
assign addr[62762]= -2067219829;
assign addr[62763]= -2045196100;
assign addr[62764]= -2020577882;
assign addr[62765]= -1993396407;
assign addr[62766]= -1963686155;
assign addr[62767]= -1931484818;
assign addr[62768]= -1896833245;
assign addr[62769]= -1859775393;
assign addr[62770]= -1820358275;
assign addr[62771]= -1778631892;
assign addr[62772]= -1734649179;
assign addr[62773]= -1688465931;
assign addr[62774]= -1640140734;
assign addr[62775]= -1589734894;
assign addr[62776]= -1537312353;
assign addr[62777]= -1482939614;
assign addr[62778]= -1426685652;
assign addr[62779]= -1368621831;
assign addr[62780]= -1308821808;
assign addr[62781]= -1247361445;
assign addr[62782]= -1184318708;
assign addr[62783]= -1119773573;
assign addr[62784]= -1053807919;
assign addr[62785]= -986505429;
assign addr[62786]= -917951481;
assign addr[62787]= -848233042;
assign addr[62788]= -777438554;
assign addr[62789]= -705657826;
assign addr[62790]= -632981917;
assign addr[62791]= -559503022;
assign addr[62792]= -485314355;
assign addr[62793]= -410510029;
assign addr[62794]= -335184940;
assign addr[62795]= -259434643;
assign addr[62796]= -183355234;
assign addr[62797]= -107043224;
assign addr[62798]= -30595422;
assign addr[62799]= 45891193;
assign addr[62800]= 122319591;
assign addr[62801]= 198592817;
assign addr[62802]= 274614114;
assign addr[62803]= 350287041;
assign addr[62804]= 425515602;
assign addr[62805]= 500204365;
assign addr[62806]= 574258580;
assign addr[62807]= 647584304;
assign addr[62808]= 720088517;
assign addr[62809]= 791679244;
assign addr[62810]= 862265664;
assign addr[62811]= 931758235;
assign addr[62812]= 1000068799;
assign addr[62813]= 1067110699;
assign addr[62814]= 1132798888;
assign addr[62815]= 1197050035;
assign addr[62816]= 1259782632;
assign addr[62817]= 1320917099;
assign addr[62818]= 1380375881;
assign addr[62819]= 1438083551;
assign addr[62820]= 1493966902;
assign addr[62821]= 1547955041;
assign addr[62822]= 1599979481;
assign addr[62823]= 1649974225;
assign addr[62824]= 1697875851;
assign addr[62825]= 1743623590;
assign addr[62826]= 1787159411;
assign addr[62827]= 1828428082;
assign addr[62828]= 1867377253;
assign addr[62829]= 1903957513;
assign addr[62830]= 1938122457;
assign addr[62831]= 1969828744;
assign addr[62832]= 1999036154;
assign addr[62833]= 2025707632;
assign addr[62834]= 2049809346;
assign addr[62835]= 2071310720;
assign addr[62836]= 2090184478;
assign addr[62837]= 2106406677;
assign addr[62838]= 2119956737;
assign addr[62839]= 2130817471;
assign addr[62840]= 2138975100;
assign addr[62841]= 2144419275;
assign addr[62842]= 2147143090;
assign addr[62843]= 2147143090;
assign addr[62844]= 2144419275;
assign addr[62845]= 2138975100;
assign addr[62846]= 2130817471;
assign addr[62847]= 2119956737;
assign addr[62848]= 2106406677;
assign addr[62849]= 2090184478;
assign addr[62850]= 2071310720;
assign addr[62851]= 2049809346;
assign addr[62852]= 2025707632;
assign addr[62853]= 1999036154;
assign addr[62854]= 1969828744;
assign addr[62855]= 1938122457;
assign addr[62856]= 1903957513;
assign addr[62857]= 1867377253;
assign addr[62858]= 1828428082;
assign addr[62859]= 1787159411;
assign addr[62860]= 1743623590;
assign addr[62861]= 1697875851;
assign addr[62862]= 1649974225;
assign addr[62863]= 1599979481;
assign addr[62864]= 1547955041;
assign addr[62865]= 1493966902;
assign addr[62866]= 1438083551;
assign addr[62867]= 1380375881;
assign addr[62868]= 1320917099;
assign addr[62869]= 1259782632;
assign addr[62870]= 1197050035;
assign addr[62871]= 1132798888;
assign addr[62872]= 1067110699;
assign addr[62873]= 1000068799;
assign addr[62874]= 931758235;
assign addr[62875]= 862265664;
assign addr[62876]= 791679244;
assign addr[62877]= 720088517;
assign addr[62878]= 647584304;
assign addr[62879]= 574258580;
assign addr[62880]= 500204365;
assign addr[62881]= 425515602;
assign addr[62882]= 350287041;
assign addr[62883]= 274614114;
assign addr[62884]= 198592817;
assign addr[62885]= 122319591;
assign addr[62886]= 45891193;
assign addr[62887]= -30595422;
assign addr[62888]= -107043224;
assign addr[62889]= -183355234;
assign addr[62890]= -259434643;
assign addr[62891]= -335184940;
assign addr[62892]= -410510029;
assign addr[62893]= -485314355;
assign addr[62894]= -559503022;
assign addr[62895]= -632981917;
assign addr[62896]= -705657826;
assign addr[62897]= -777438554;
assign addr[62898]= -848233042;
assign addr[62899]= -917951481;
assign addr[62900]= -986505429;
assign addr[62901]= -1053807919;
assign addr[62902]= -1119773573;
assign addr[62903]= -1184318708;
assign addr[62904]= -1247361445;
assign addr[62905]= -1308821808;
assign addr[62906]= -1368621831;
assign addr[62907]= -1426685652;
assign addr[62908]= -1482939614;
assign addr[62909]= -1537312353;
assign addr[62910]= -1589734894;
assign addr[62911]= -1640140734;
assign addr[62912]= -1688465931;
assign addr[62913]= -1734649179;
assign addr[62914]= -1778631892;
assign addr[62915]= -1820358275;
assign addr[62916]= -1859775393;
assign addr[62917]= -1896833245;
assign addr[62918]= -1931484818;
assign addr[62919]= -1963686155;
assign addr[62920]= -1993396407;
assign addr[62921]= -2020577882;
assign addr[62922]= -2045196100;
assign addr[62923]= -2067219829;
assign addr[62924]= -2086621133;
assign addr[62925]= -2103375398;
assign addr[62926]= -2117461370;
assign addr[62927]= -2128861181;
assign addr[62928]= -2137560369;
assign addr[62929]= -2143547897;
assign addr[62930]= -2146816171;
assign addr[62931]= -2147361045;
assign addr[62932]= -2145181827;
assign addr[62933]= -2140281282;
assign addr[62934]= -2132665626;
assign addr[62935]= -2122344521;
assign addr[62936]= -2109331059;
assign addr[62937]= -2093641749;
assign addr[62938]= -2075296495;
assign addr[62939]= -2054318569;
assign addr[62940]= -2030734582;
assign addr[62941]= -2004574453;
assign addr[62942]= -1975871368;
assign addr[62943]= -1944661739;
assign addr[62944]= -1910985158;
assign addr[62945]= -1874884346;
assign addr[62946]= -1836405100;
assign addr[62947]= -1795596234;
assign addr[62948]= -1752509516;
assign addr[62949]= -1707199606;
assign addr[62950]= -1659723983;
assign addr[62951]= -1610142873;
assign addr[62952]= -1558519173;
assign addr[62953]= -1504918373;
assign addr[62954]= -1449408469;
assign addr[62955]= -1392059879;
assign addr[62956]= -1332945355;
assign addr[62957]= -1272139887;
assign addr[62958]= -1209720613;
assign addr[62959]= -1145766716;
assign addr[62960]= -1080359326;
assign addr[62961]= -1013581418;
assign addr[62962]= -945517704;
assign addr[62963]= -876254528;
assign addr[62964]= -805879757;
assign addr[62965]= -734482665;
assign addr[62966]= -662153826;
assign addr[62967]= -588984994;
assign addr[62968]= -515068990;
assign addr[62969]= -440499581;
assign addr[62970]= -365371365;
assign addr[62971]= -289779648;
assign addr[62972]= -213820322;
assign addr[62973]= -137589750;
assign addr[62974]= -61184634;
assign addr[62975]= 15298099;
assign addr[62976]= 91761426;
assign addr[62977]= 168108346;
assign addr[62978]= 244242007;
assign addr[62979]= 320065829;
assign addr[62980]= 395483624;
assign addr[62981]= 470399716;
assign addr[62982]= 544719071;
assign addr[62983]= 618347408;
assign addr[62984]= 691191324;
assign addr[62985]= 763158411;
assign addr[62986]= 834157373;
assign addr[62987]= 904098143;
assign addr[62988]= 972891995;
assign addr[62989]= 1040451659;
assign addr[62990]= 1106691431;
assign addr[62991]= 1171527280;
assign addr[62992]= 1234876957;
assign addr[62993]= 1296660098;
assign addr[62994]= 1356798326;
assign addr[62995]= 1415215352;
assign addr[62996]= 1471837070;
assign addr[62997]= 1526591649;
assign addr[62998]= 1579409630;
assign addr[62999]= 1630224009;
assign addr[63000]= 1678970324;
assign addr[63001]= 1725586737;
assign addr[63002]= 1770014111;
assign addr[63003]= 1812196087;
assign addr[63004]= 1852079154;
assign addr[63005]= 1889612716;
assign addr[63006]= 1924749160;
assign addr[63007]= 1957443913;
assign addr[63008]= 1987655498;
assign addr[63009]= 2015345591;
assign addr[63010]= 2040479063;
assign addr[63011]= 2063024031;
assign addr[63012]= 2082951896;
assign addr[63013]= 2100237377;
assign addr[63014]= 2114858546;
assign addr[63015]= 2126796855;
assign addr[63016]= 2136037160;
assign addr[63017]= 2142567738;
assign addr[63018]= 2146380306;
assign addr[63019]= 2147470025;
assign addr[63020]= 2145835515;
assign addr[63021]= 2141478848;
assign addr[63022]= 2134405552;
assign addr[63023]= 2124624598;
assign addr[63024]= 2112148396;
assign addr[63025]= 2096992772;
assign addr[63026]= 2079176953;
assign addr[63027]= 2058723538;
assign addr[63028]= 2035658475;
assign addr[63029]= 2010011024;
assign addr[63030]= 1981813720;
assign addr[63031]= 1951102334;
assign addr[63032]= 1917915825;
assign addr[63033]= 1882296293;
assign addr[63034]= 1844288924;
assign addr[63035]= 1803941934;
assign addr[63036]= 1761306505;
assign addr[63037]= 1716436725;
assign addr[63038]= 1669389513;
assign addr[63039]= 1620224553;
assign addr[63040]= 1569004214;
assign addr[63041]= 1515793473;
assign addr[63042]= 1460659832;
assign addr[63043]= 1403673233;
assign addr[63044]= 1344905966;
assign addr[63045]= 1284432584;
assign addr[63046]= 1222329801;
assign addr[63047]= 1158676398;
assign addr[63048]= 1093553126;
assign addr[63049]= 1027042599;
assign addr[63050]= 959229189;
assign addr[63051]= 890198924;
assign addr[63052]= 820039373;
assign addr[63053]= 748839539;
assign addr[63054]= 676689746;
assign addr[63055]= 603681519;
assign addr[63056]= 529907477;
assign addr[63057]= 455461206;
assign addr[63058]= 380437148;
assign addr[63059]= 304930476;
assign addr[63060]= 229036977;
assign addr[63061]= 152852926;
assign addr[63062]= 76474970;
assign addr[63063]= 0;
assign addr[63064]= -76474970;
assign addr[63065]= -152852926;
assign addr[63066]= -229036977;
assign addr[63067]= -304930476;
assign addr[63068]= -380437148;
assign addr[63069]= -455461206;
assign addr[63070]= -529907477;
assign addr[63071]= -603681519;
assign addr[63072]= -676689746;
assign addr[63073]= -748839539;
assign addr[63074]= -820039373;
assign addr[63075]= -890198924;
assign addr[63076]= -959229189;
assign addr[63077]= -1027042599;
assign addr[63078]= -1093553126;
assign addr[63079]= -1158676398;
assign addr[63080]= -1222329801;
assign addr[63081]= -1284432584;
assign addr[63082]= -1344905966;
assign addr[63083]= -1403673233;
assign addr[63084]= -1460659832;
assign addr[63085]= -1515793473;
assign addr[63086]= -1569004214;
assign addr[63087]= -1620224553;
assign addr[63088]= -1669389513;
assign addr[63089]= -1716436725;
assign addr[63090]= -1761306505;
assign addr[63091]= -1803941934;
assign addr[63092]= -1844288924;
assign addr[63093]= -1882296293;
assign addr[63094]= -1917915825;
assign addr[63095]= -1951102334;
assign addr[63096]= -1981813720;
assign addr[63097]= -2010011024;
assign addr[63098]= -2035658475;
assign addr[63099]= -2058723538;
assign addr[63100]= -2079176953;
assign addr[63101]= -2096992772;
assign addr[63102]= -2112148396;
assign addr[63103]= -2124624598;
assign addr[63104]= -2134405552;
assign addr[63105]= -2141478848;
assign addr[63106]= -2145835515;
assign addr[63107]= -2147470025;
assign addr[63108]= -2146380306;
assign addr[63109]= -2142567738;
assign addr[63110]= -2136037160;
assign addr[63111]= -2126796855;
assign addr[63112]= -2114858546;
assign addr[63113]= -2100237377;
assign addr[63114]= -2082951896;
assign addr[63115]= -2063024031;
assign addr[63116]= -2040479063;
assign addr[63117]= -2015345591;
assign addr[63118]= -1987655498;
assign addr[63119]= -1957443913;
assign addr[63120]= -1924749160;
assign addr[63121]= -1889612716;
assign addr[63122]= -1852079154;
assign addr[63123]= -1812196087;
assign addr[63124]= -1770014111;
assign addr[63125]= -1725586737;
assign addr[63126]= -1678970324;
assign addr[63127]= -1630224009;
assign addr[63128]= -1579409630;
assign addr[63129]= -1526591649;
assign addr[63130]= -1471837070;
assign addr[63131]= -1415215352;
assign addr[63132]= -1356798326;
assign addr[63133]= -1296660098;
assign addr[63134]= -1234876957;
assign addr[63135]= -1171527280;
assign addr[63136]= -1106691431;
assign addr[63137]= -1040451659;
assign addr[63138]= -972891995;
assign addr[63139]= -904098143;
assign addr[63140]= -834157373;
assign addr[63141]= -763158411;
assign addr[63142]= -691191324;
assign addr[63143]= -618347408;
assign addr[63144]= -544719071;
assign addr[63145]= -470399716;
assign addr[63146]= -395483624;
assign addr[63147]= -320065829;
assign addr[63148]= -244242007;
assign addr[63149]= -168108346;
assign addr[63150]= -91761426;
assign addr[63151]= -15298099;
assign addr[63152]= 61184634;
assign addr[63153]= 137589750;
assign addr[63154]= 213820322;
assign addr[63155]= 289779648;
assign addr[63156]= 365371365;
assign addr[63157]= 440499581;
assign addr[63158]= 515068990;
assign addr[63159]= 588984994;
assign addr[63160]= 662153826;
assign addr[63161]= 734482665;
assign addr[63162]= 805879757;
assign addr[63163]= 876254528;
assign addr[63164]= 945517704;
assign addr[63165]= 1013581418;
assign addr[63166]= 1080359326;
assign addr[63167]= 1145766716;
assign addr[63168]= 1209720613;
assign addr[63169]= 1272139887;
assign addr[63170]= 1332945355;
assign addr[63171]= 1392059879;
assign addr[63172]= 1449408469;
assign addr[63173]= 1504918373;
assign addr[63174]= 1558519173;
assign addr[63175]= 1610142873;
assign addr[63176]= 1659723983;
assign addr[63177]= 1707199606;
assign addr[63178]= 1752509516;
assign addr[63179]= 1795596234;
assign addr[63180]= 1836405100;
assign addr[63181]= 1874884346;
assign addr[63182]= 1910985158;
assign addr[63183]= 1944661739;
assign addr[63184]= 1975871368;
assign addr[63185]= 2004574453;
assign addr[63186]= 2030734582;
assign addr[63187]= 2054318569;
assign addr[63188]= 2075296495;
assign addr[63189]= 2093641749;
assign addr[63190]= 2109331059;
assign addr[63191]= 2122344521;
assign addr[63192]= 2132665626;
assign addr[63193]= 2140281282;
assign addr[63194]= 2145181827;
assign addr[63195]= 2147361045;
assign addr[63196]= 2146816171;
assign addr[63197]= 2143547897;
assign addr[63198]= 2137560369;
assign addr[63199]= 2128861181;
assign addr[63200]= 2117461370;
assign addr[63201]= 2103375398;
assign addr[63202]= 2086621133;
assign addr[63203]= 2067219829;
assign addr[63204]= 2045196100;
assign addr[63205]= 2020577882;
assign addr[63206]= 1993396407;
assign addr[63207]= 1963686155;
assign addr[63208]= 1931484818;
assign addr[63209]= 1896833245;
assign addr[63210]= 1859775393;
assign addr[63211]= 1820358275;
assign addr[63212]= 1778631892;
assign addr[63213]= 1734649179;
assign addr[63214]= 1688465931;
assign addr[63215]= 1640140734;
assign addr[63216]= 1589734894;
assign addr[63217]= 1537312353;
assign addr[63218]= 1482939614;
assign addr[63219]= 1426685652;
assign addr[63220]= 1368621831;
assign addr[63221]= 1308821808;
assign addr[63222]= 1247361445;
assign addr[63223]= 1184318708;
assign addr[63224]= 1119773573;
assign addr[63225]= 1053807919;
assign addr[63226]= 986505429;
assign addr[63227]= 917951481;
assign addr[63228]= 848233042;
assign addr[63229]= 777438554;
assign addr[63230]= 705657826;
assign addr[63231]= 632981917;
assign addr[63232]= 559503022;
assign addr[63233]= 485314355;
assign addr[63234]= 410510029;
assign addr[63235]= 335184940;
assign addr[63236]= 259434643;
assign addr[63237]= 183355234;
assign addr[63238]= 107043224;
assign addr[63239]= 30595422;
assign addr[63240]= -45891193;
assign addr[63241]= -122319591;
assign addr[63242]= -198592817;
assign addr[63243]= -274614114;
assign addr[63244]= -350287041;
assign addr[63245]= -425515602;
assign addr[63246]= -500204365;
assign addr[63247]= -574258580;
assign addr[63248]= -647584304;
assign addr[63249]= -720088517;
assign addr[63250]= -791679244;
assign addr[63251]= -862265664;
assign addr[63252]= -931758235;
assign addr[63253]= -1000068799;
assign addr[63254]= -1067110699;
assign addr[63255]= -1132798888;
assign addr[63256]= -1197050035;
assign addr[63257]= -1259782632;
assign addr[63258]= -1320917099;
assign addr[63259]= -1380375881;
assign addr[63260]= -1438083551;
assign addr[63261]= -1493966902;
assign addr[63262]= -1547955041;
assign addr[63263]= -1599979481;
assign addr[63264]= -1649974225;
assign addr[63265]= -1697875851;
assign addr[63266]= -1743623590;
assign addr[63267]= -1787159411;
assign addr[63268]= -1828428082;
assign addr[63269]= -1867377253;
assign addr[63270]= -1903957513;
assign addr[63271]= -1938122457;
assign addr[63272]= -1969828744;
assign addr[63273]= -1999036154;
assign addr[63274]= -2025707632;
assign addr[63275]= -2049809346;
assign addr[63276]= -2071310720;
assign addr[63277]= -2090184478;
assign addr[63278]= -2106406677;
assign addr[63279]= -2119956737;
assign addr[63280]= -2130817471;
assign addr[63281]= -2138975100;
assign addr[63282]= -2144419275;
assign addr[63283]= -2147143090;
assign addr[63284]= -2147143090;
assign addr[63285]= -2144419275;
assign addr[63286]= -2138975100;
assign addr[63287]= -2130817471;
assign addr[63288]= -2119956737;
assign addr[63289]= -2106406677;
assign addr[63290]= -2090184478;
assign addr[63291]= -2071310720;
assign addr[63292]= -2049809346;
assign addr[63293]= -2025707632;
assign addr[63294]= -1999036154;
assign addr[63295]= -1969828744;
assign addr[63296]= -1938122457;
assign addr[63297]= -1903957513;
assign addr[63298]= -1867377253;
assign addr[63299]= -1828428082;
assign addr[63300]= -1787159411;
assign addr[63301]= -1743623590;
assign addr[63302]= -1697875851;
assign addr[63303]= -1649974225;
assign addr[63304]= -1599979481;
assign addr[63305]= -1547955041;
assign addr[63306]= -1493966902;
assign addr[63307]= -1438083551;
assign addr[63308]= -1380375881;
assign addr[63309]= -1320917099;
assign addr[63310]= -1259782632;
assign addr[63311]= -1197050035;
assign addr[63312]= -1132798888;
assign addr[63313]= -1067110699;
assign addr[63314]= -1000068799;
assign addr[63315]= -931758235;
assign addr[63316]= -862265664;
assign addr[63317]= -791679244;
assign addr[63318]= -720088517;
assign addr[63319]= -647584304;
assign addr[63320]= -574258580;
assign addr[63321]= -500204365;
assign addr[63322]= -425515602;
assign addr[63323]= -350287041;
assign addr[63324]= -274614114;
assign addr[63325]= -198592817;
assign addr[63326]= -122319591;
assign addr[63327]= -45891193;
assign addr[63328]= 30595422;
assign addr[63329]= 107043224;
assign addr[63330]= 183355234;
assign addr[63331]= 259434643;
assign addr[63332]= 335184940;
assign addr[63333]= 410510029;
assign addr[63334]= 485314355;
assign addr[63335]= 559503022;
assign addr[63336]= 632981917;
assign addr[63337]= 705657826;
assign addr[63338]= 777438554;
assign addr[63339]= 848233042;
assign addr[63340]= 917951481;
assign addr[63341]= 986505429;
assign addr[63342]= 1053807919;
assign addr[63343]= 1119773573;
assign addr[63344]= 1184318708;
assign addr[63345]= 1247361445;
assign addr[63346]= 1308821808;
assign addr[63347]= 1368621831;
assign addr[63348]= 1426685652;
assign addr[63349]= 1482939614;
assign addr[63350]= 1537312353;
assign addr[63351]= 1589734894;
assign addr[63352]= 1640140734;
assign addr[63353]= 1688465931;
assign addr[63354]= 1734649179;
assign addr[63355]= 1778631892;
assign addr[63356]= 1820358275;
assign addr[63357]= 1859775393;
assign addr[63358]= 1896833245;
assign addr[63359]= 1931484818;
assign addr[63360]= 1963686155;
assign addr[63361]= 1993396407;
assign addr[63362]= 2020577882;
assign addr[63363]= 2045196100;
assign addr[63364]= 2067219829;
assign addr[63365]= 2086621133;
assign addr[63366]= 2103375398;
assign addr[63367]= 2117461370;
assign addr[63368]= 2128861181;
assign addr[63369]= 2137560369;
assign addr[63370]= 2143547897;
assign addr[63371]= 2146816171;
assign addr[63372]= 2147361045;
assign addr[63373]= 2145181827;
assign addr[63374]= 2140281282;
assign addr[63375]= 2132665626;
assign addr[63376]= 2122344521;
assign addr[63377]= 2109331059;
assign addr[63378]= 2093641749;
assign addr[63379]= 2075296495;
assign addr[63380]= 2054318569;
assign addr[63381]= 2030734582;
assign addr[63382]= 2004574453;
assign addr[63383]= 1975871368;
assign addr[63384]= 1944661739;
assign addr[63385]= 1910985158;
assign addr[63386]= 1874884346;
assign addr[63387]= 1836405100;
assign addr[63388]= 1795596234;
assign addr[63389]= 1752509516;
assign addr[63390]= 1707199606;
assign addr[63391]= 1659723983;
assign addr[63392]= 1610142873;
assign addr[63393]= 1558519173;
assign addr[63394]= 1504918373;
assign addr[63395]= 1449408469;
assign addr[63396]= 1392059879;
assign addr[63397]= 1332945355;
assign addr[63398]= 1272139887;
assign addr[63399]= 1209720613;
assign addr[63400]= 1145766716;
assign addr[63401]= 1080359326;
assign addr[63402]= 1013581418;
assign addr[63403]= 945517704;
assign addr[63404]= 876254528;
assign addr[63405]= 805879757;
assign addr[63406]= 734482665;
assign addr[63407]= 662153826;
assign addr[63408]= 588984994;
assign addr[63409]= 515068990;
assign addr[63410]= 440499581;
assign addr[63411]= 365371365;
assign addr[63412]= 289779648;
assign addr[63413]= 213820322;
assign addr[63414]= 137589750;
assign addr[63415]= 61184634;
assign addr[63416]= -15298099;
assign addr[63417]= -91761426;
assign addr[63418]= -168108346;
assign addr[63419]= -244242007;
assign addr[63420]= -320065829;
assign addr[63421]= -395483624;
assign addr[63422]= -470399716;
assign addr[63423]= -544719071;
assign addr[63424]= -618347408;
assign addr[63425]= -691191324;
assign addr[63426]= -763158411;
assign addr[63427]= -834157373;
assign addr[63428]= -904098143;
assign addr[63429]= -972891995;
assign addr[63430]= -1040451659;
assign addr[63431]= -1106691431;
assign addr[63432]= -1171527280;
assign addr[63433]= -1234876957;
assign addr[63434]= -1296660098;
assign addr[63435]= -1356798326;
assign addr[63436]= -1415215352;
assign addr[63437]= -1471837070;
assign addr[63438]= -1526591649;
assign addr[63439]= -1579409630;
assign addr[63440]= -1630224009;
assign addr[63441]= -1678970324;
assign addr[63442]= -1725586737;
assign addr[63443]= -1770014111;
assign addr[63444]= -1812196087;
assign addr[63445]= -1852079154;
assign addr[63446]= -1889612716;
assign addr[63447]= -1924749160;
assign addr[63448]= -1957443913;
assign addr[63449]= -1987655498;
assign addr[63450]= -2015345591;
assign addr[63451]= -2040479063;
assign addr[63452]= -2063024031;
assign addr[63453]= -2082951896;
assign addr[63454]= -2100237377;
assign addr[63455]= -2114858546;
assign addr[63456]= -2126796855;
assign addr[63457]= -2136037160;
assign addr[63458]= -2142567738;
assign addr[63459]= -2146380306;
assign addr[63460]= -2147470025;
assign addr[63461]= -2145835515;
assign addr[63462]= -2141478848;
assign addr[63463]= -2134405552;
assign addr[63464]= -2124624598;
assign addr[63465]= -2112148396;
assign addr[63466]= -2096992772;
assign addr[63467]= -2079176953;
assign addr[63468]= -2058723538;
assign addr[63469]= -2035658475;
assign addr[63470]= -2010011024;
assign addr[63471]= -1981813720;
assign addr[63472]= -1951102334;
assign addr[63473]= -1917915825;
assign addr[63474]= -1882296293;
assign addr[63475]= -1844288924;
assign addr[63476]= -1803941934;
assign addr[63477]= -1761306505;
assign addr[63478]= -1716436725;
assign addr[63479]= -1669389513;
assign addr[63480]= -1620224553;
assign addr[63481]= -1569004214;
assign addr[63482]= -1515793473;
assign addr[63483]= -1460659832;
assign addr[63484]= -1403673233;
assign addr[63485]= -1344905966;
assign addr[63486]= -1284432584;
assign addr[63487]= -1222329801;
assign addr[63488]= -1158676398;
assign addr[63489]= -1093553126;
assign addr[63490]= -1027042599;
assign addr[63491]= -959229189;
assign addr[63492]= -890198924;
assign addr[63493]= -820039373;
assign addr[63494]= -748839539;
assign addr[63495]= -676689746;
assign addr[63496]= -603681519;
assign addr[63497]= -529907477;
assign addr[63498]= -455461206;
assign addr[63499]= -380437148;
assign addr[63500]= -304930476;
assign addr[63501]= -229036977;
assign addr[63502]= -152852926;
assign addr[63503]= -76474970;
assign addr[63504]= 0;
assign addr[63505]= 76474970;
assign addr[63506]= 152852926;
assign addr[63507]= 229036977;
assign addr[63508]= 304930476;
assign addr[63509]= 380437148;
assign addr[63510]= 455461206;
assign addr[63511]= 529907477;
assign addr[63512]= 603681519;
assign addr[63513]= 676689746;
assign addr[63514]= 748839539;
assign addr[63515]= 820039373;
assign addr[63516]= 890198924;
assign addr[63517]= 959229189;
assign addr[63518]= 1027042599;
assign addr[63519]= 1093553126;
assign addr[63520]= 1158676398;
assign addr[63521]= 1222329801;
assign addr[63522]= 1284432584;
assign addr[63523]= 1344905966;
assign addr[63524]= 1403673233;
assign addr[63525]= 1460659832;
assign addr[63526]= 1515793473;
assign addr[63527]= 1569004214;
assign addr[63528]= 1620224553;
assign addr[63529]= 1669389513;
assign addr[63530]= 1716436725;
assign addr[63531]= 1761306505;
assign addr[63532]= 1803941934;
assign addr[63533]= 1844288924;
assign addr[63534]= 1882296293;
assign addr[63535]= 1917915825;
assign addr[63536]= 1951102334;
assign addr[63537]= 1981813720;
assign addr[63538]= 2010011024;
assign addr[63539]= 2035658475;
assign addr[63540]= 2058723538;
assign addr[63541]= 2079176953;
assign addr[63542]= 2096992772;
assign addr[63543]= 2112148396;
assign addr[63544]= 2124624598;
assign addr[63545]= 2134405552;
assign addr[63546]= 2141478848;
assign addr[63547]= 2145835515;
assign addr[63548]= 2147470025;
assign addr[63549]= 2146380306;
assign addr[63550]= 2142567738;
assign addr[63551]= 2136037160;
assign addr[63552]= 2126796855;
assign addr[63553]= 2114858546;
assign addr[63554]= 2100237377;
assign addr[63555]= 2082951896;
assign addr[63556]= 2063024031;
assign addr[63557]= 2040479063;
assign addr[63558]= 2015345591;
assign addr[63559]= 1987655498;
assign addr[63560]= 1957443913;
assign addr[63561]= 1924749160;
assign addr[63562]= 1889612716;
assign addr[63563]= 1852079154;
assign addr[63564]= 1812196087;
assign addr[63565]= 1770014111;
assign addr[63566]= 1725586737;
assign addr[63567]= 1678970324;
assign addr[63568]= 1630224009;
assign addr[63569]= 1579409630;
assign addr[63570]= 1526591649;
assign addr[63571]= 1471837070;
assign addr[63572]= 1415215352;
assign addr[63573]= 1356798326;
assign addr[63574]= 1296660098;
assign addr[63575]= 1234876957;
assign addr[63576]= 1171527280;
assign addr[63577]= 1106691431;
assign addr[63578]= 1040451659;
assign addr[63579]= 972891995;
assign addr[63580]= 904098143;
assign addr[63581]= 834157373;
assign addr[63582]= 763158411;
assign addr[63583]= 691191324;
assign addr[63584]= 618347408;
assign addr[63585]= 544719071;
assign addr[63586]= 470399716;
assign addr[63587]= 395483624;
assign addr[63588]= 320065829;
assign addr[63589]= 244242007;
assign addr[63590]= 168108346;
assign addr[63591]= 91761426;
assign addr[63592]= 15298099;
assign addr[63593]= -61184634;
assign addr[63594]= -137589750;
assign addr[63595]= -213820322;
assign addr[63596]= -289779648;
assign addr[63597]= -365371365;
assign addr[63598]= -440499581;
assign addr[63599]= -515068990;
assign addr[63600]= -588984994;
assign addr[63601]= -662153826;
assign addr[63602]= -734482665;
assign addr[63603]= -805879757;
assign addr[63604]= -876254528;
assign addr[63605]= -945517704;
assign addr[63606]= -1013581418;
assign addr[63607]= -1080359326;
assign addr[63608]= -1145766716;
assign addr[63609]= -1209720613;
assign addr[63610]= -1272139887;
assign addr[63611]= -1332945355;
assign addr[63612]= -1392059879;
assign addr[63613]= -1449408469;
assign addr[63614]= -1504918373;
assign addr[63615]= -1558519173;
assign addr[63616]= -1610142873;
assign addr[63617]= -1659723983;
assign addr[63618]= -1707199606;
assign addr[63619]= -1752509516;
assign addr[63620]= -1795596234;
assign addr[63621]= -1836405100;
assign addr[63622]= -1874884346;
assign addr[63623]= -1910985158;
assign addr[63624]= -1944661739;
assign addr[63625]= -1975871368;
assign addr[63626]= -2004574453;
assign addr[63627]= -2030734582;
assign addr[63628]= -2054318569;
assign addr[63629]= -2075296495;
assign addr[63630]= -2093641749;
assign addr[63631]= -2109331059;
assign addr[63632]= -2122344521;
assign addr[63633]= -2132665626;
assign addr[63634]= -2140281282;
assign addr[63635]= -2145181827;
assign addr[63636]= -2147361045;
assign addr[63637]= -2146816171;
assign addr[63638]= -2143547897;
assign addr[63639]= -2137560369;
assign addr[63640]= -2128861181;
assign addr[63641]= -2117461370;
assign addr[63642]= -2103375398;
assign addr[63643]= -2086621133;
assign addr[63644]= -2067219829;
assign addr[63645]= -2045196100;
assign addr[63646]= -2020577882;
assign addr[63647]= -1993396407;
assign addr[63648]= -1963686155;
assign addr[63649]= -1931484818;
assign addr[63650]= -1896833245;
assign addr[63651]= -1859775393;
assign addr[63652]= -1820358275;
assign addr[63653]= -1778631892;
assign addr[63654]= -1734649179;
assign addr[63655]= -1688465931;
assign addr[63656]= -1640140734;
assign addr[63657]= -1589734894;
assign addr[63658]= -1537312353;
assign addr[63659]= -1482939614;
assign addr[63660]= -1426685652;
assign addr[63661]= -1368621831;
assign addr[63662]= -1308821808;
assign addr[63663]= -1247361445;
assign addr[63664]= -1184318708;
assign addr[63665]= -1119773573;
assign addr[63666]= -1053807919;
assign addr[63667]= -986505429;
assign addr[63668]= -917951481;
assign addr[63669]= -848233042;
assign addr[63670]= -777438554;
assign addr[63671]= -705657826;
assign addr[63672]= -632981917;
assign addr[63673]= -559503022;
assign addr[63674]= -485314355;
assign addr[63675]= -410510029;
assign addr[63676]= -335184940;
assign addr[63677]= -259434643;
assign addr[63678]= -183355234;
assign addr[63679]= -107043224;
assign addr[63680]= -30595422;
assign addr[63681]= 45891193;
assign addr[63682]= 122319591;
assign addr[63683]= 198592817;
assign addr[63684]= 274614114;
assign addr[63685]= 350287041;
assign addr[63686]= 425515602;
assign addr[63687]= 500204365;
assign addr[63688]= 574258580;
assign addr[63689]= 647584304;
assign addr[63690]= 720088517;
assign addr[63691]= 791679244;
assign addr[63692]= 862265664;
assign addr[63693]= 931758235;
assign addr[63694]= 1000068799;
assign addr[63695]= 1067110699;
assign addr[63696]= 1132798888;
assign addr[63697]= 1197050035;
assign addr[63698]= 1259782632;
assign addr[63699]= 1320917099;
assign addr[63700]= 1380375881;
assign addr[63701]= 1438083551;
assign addr[63702]= 1493966902;
assign addr[63703]= 1547955041;
assign addr[63704]= 1599979481;
assign addr[63705]= 1649974225;
assign addr[63706]= 1697875851;
assign addr[63707]= 1743623590;
assign addr[63708]= 1787159411;
assign addr[63709]= 1828428082;
assign addr[63710]= 1867377253;
assign addr[63711]= 1903957513;
assign addr[63712]= 1938122457;
assign addr[63713]= 1969828744;
assign addr[63714]= 1999036154;
assign addr[63715]= 2025707632;
assign addr[63716]= 2049809346;
assign addr[63717]= 2071310720;
assign addr[63718]= 2090184478;
assign addr[63719]= 2106406677;
assign addr[63720]= 2119956737;
assign addr[63721]= 2130817471;
assign addr[63722]= 2138975100;
assign addr[63723]= 2144419275;
assign addr[63724]= 2147143090;
assign addr[63725]= 2147143090;
assign addr[63726]= 2144419275;
assign addr[63727]= 2138975100;
assign addr[63728]= 2130817471;
assign addr[63729]= 2119956737;
assign addr[63730]= 2106406677;
assign addr[63731]= 2090184478;
assign addr[63732]= 2071310720;
assign addr[63733]= 2049809346;
assign addr[63734]= 2025707632;
assign addr[63735]= 1999036154;
assign addr[63736]= 1969828744;
assign addr[63737]= 1938122457;
assign addr[63738]= 1903957513;
assign addr[63739]= 1867377253;
assign addr[63740]= 1828428082;
assign addr[63741]= 1787159411;
assign addr[63742]= 1743623590;
assign addr[63743]= 1697875851;
assign addr[63744]= 1649974225;
assign addr[63745]= 1599979481;
assign addr[63746]= 1547955041;
assign addr[63747]= 1493966902;
assign addr[63748]= 1438083551;
assign addr[63749]= 1380375881;
assign addr[63750]= 1320917099;
assign addr[63751]= 1259782632;
assign addr[63752]= 1197050035;
assign addr[63753]= 1132798888;
assign addr[63754]= 1067110699;
assign addr[63755]= 1000068799;
assign addr[63756]= 931758235;
assign addr[63757]= 862265664;
assign addr[63758]= 791679244;
assign addr[63759]= 720088517;
assign addr[63760]= 647584304;
assign addr[63761]= 574258580;
assign addr[63762]= 500204365;
assign addr[63763]= 425515602;
assign addr[63764]= 350287041;
assign addr[63765]= 274614114;
assign addr[63766]= 198592817;
assign addr[63767]= 122319591;
assign addr[63768]= 45891193;
assign addr[63769]= -30595422;
assign addr[63770]= -107043224;
assign addr[63771]= -183355234;
assign addr[63772]= -259434643;
assign addr[63773]= -335184940;
assign addr[63774]= -410510029;
assign addr[63775]= -485314355;
assign addr[63776]= -559503022;
assign addr[63777]= -632981917;
assign addr[63778]= -705657826;
assign addr[63779]= -777438554;
assign addr[63780]= -848233042;
assign addr[63781]= -917951481;
assign addr[63782]= -986505429;
assign addr[63783]= -1053807919;
assign addr[63784]= -1119773573;
assign addr[63785]= -1184318708;
assign addr[63786]= -1247361445;
assign addr[63787]= -1308821808;
assign addr[63788]= -1368621831;
assign addr[63789]= -1426685652;
assign addr[63790]= -1482939614;
assign addr[63791]= -1537312353;
assign addr[63792]= -1589734894;
assign addr[63793]= -1640140734;
assign addr[63794]= -1688465931;
assign addr[63795]= -1734649179;
assign addr[63796]= -1778631892;
assign addr[63797]= -1820358275;
assign addr[63798]= -1859775393;
assign addr[63799]= -1896833245;
assign addr[63800]= -1931484818;
assign addr[63801]= -1963686155;
assign addr[63802]= -1993396407;
assign addr[63803]= -2020577882;
assign addr[63804]= -2045196100;
assign addr[63805]= -2067219829;
assign addr[63806]= -2086621133;
assign addr[63807]= -2103375398;
assign addr[63808]= -2117461370;
assign addr[63809]= -2128861181;
assign addr[63810]= -2137560369;
assign addr[63811]= -2143547897;
assign addr[63812]= -2146816171;
assign addr[63813]= -2147361045;
assign addr[63814]= -2145181827;
assign addr[63815]= -2140281282;
assign addr[63816]= -2132665626;
assign addr[63817]= -2122344521;
assign addr[63818]= -2109331059;
assign addr[63819]= -2093641749;
assign addr[63820]= -2075296495;
assign addr[63821]= -2054318569;
assign addr[63822]= -2030734582;
assign addr[63823]= -2004574453;
assign addr[63824]= -1975871368;
assign addr[63825]= -1944661739;
assign addr[63826]= -1910985158;
assign addr[63827]= -1874884346;
assign addr[63828]= -1836405100;
assign addr[63829]= -1795596234;
assign addr[63830]= -1752509516;
assign addr[63831]= -1707199606;
assign addr[63832]= -1659723983;
assign addr[63833]= -1610142873;
assign addr[63834]= -1558519173;
assign addr[63835]= -1504918373;
assign addr[63836]= -1449408469;
assign addr[63837]= -1392059879;
assign addr[63838]= -1332945355;
assign addr[63839]= -1272139887;
assign addr[63840]= -1209720613;
assign addr[63841]= -1145766716;
assign addr[63842]= -1080359326;
assign addr[63843]= -1013581418;
assign addr[63844]= -945517704;
assign addr[63845]= -876254528;
assign addr[63846]= -805879757;
assign addr[63847]= -734482665;
assign addr[63848]= -662153826;
assign addr[63849]= -588984994;
assign addr[63850]= -515068990;
assign addr[63851]= -440499581;
assign addr[63852]= -365371365;
assign addr[63853]= -289779648;
assign addr[63854]= -213820322;
assign addr[63855]= -137589750;
assign addr[63856]= -61184634;
assign addr[63857]= 15298099;
assign addr[63858]= 91761426;
assign addr[63859]= 168108346;
assign addr[63860]= 244242007;
assign addr[63861]= 320065829;
assign addr[63862]= 395483624;
assign addr[63863]= 470399716;
assign addr[63864]= 544719071;
assign addr[63865]= 618347408;
assign addr[63866]= 691191324;
assign addr[63867]= 763158411;
assign addr[63868]= 834157373;
assign addr[63869]= 904098143;
assign addr[63870]= 972891995;
assign addr[63871]= 1040451659;
assign addr[63872]= 1106691431;
assign addr[63873]= 1171527280;
assign addr[63874]= 1234876957;
assign addr[63875]= 1296660098;
assign addr[63876]= 1356798326;
assign addr[63877]= 1415215352;
assign addr[63878]= 1471837070;
assign addr[63879]= 1526591649;
assign addr[63880]= 1579409630;
assign addr[63881]= 1630224009;
assign addr[63882]= 1678970324;
assign addr[63883]= 1725586737;
assign addr[63884]= 1770014111;
assign addr[63885]= 1812196087;
assign addr[63886]= 1852079154;
assign addr[63887]= 1889612716;
assign addr[63888]= 1924749160;
assign addr[63889]= 1957443913;
assign addr[63890]= 1987655498;
assign addr[63891]= 2015345591;
assign addr[63892]= 2040479063;
assign addr[63893]= 2063024031;
assign addr[63894]= 2082951896;
assign addr[63895]= 2100237377;
assign addr[63896]= 2114858546;
assign addr[63897]= 2126796855;
assign addr[63898]= 2136037160;
assign addr[63899]= 2142567738;
assign addr[63900]= 2146380306;
assign addr[63901]= 2147470025;
assign addr[63902]= 2145835515;
assign addr[63903]= 2141478848;
assign addr[63904]= 2134405552;
assign addr[63905]= 2124624598;
assign addr[63906]= 2112148396;
assign addr[63907]= 2096992772;
assign addr[63908]= 2079176953;
assign addr[63909]= 2058723538;
assign addr[63910]= 2035658475;
assign addr[63911]= 2010011024;
assign addr[63912]= 1981813720;
assign addr[63913]= 1951102334;
assign addr[63914]= 1917915825;
assign addr[63915]= 1882296293;
assign addr[63916]= 1844288924;
assign addr[63917]= 1803941934;
assign addr[63918]= 1761306505;
assign addr[63919]= 1716436725;
assign addr[63920]= 1669389513;
assign addr[63921]= 1620224553;
assign addr[63922]= 1569004214;
assign addr[63923]= 1515793473;
assign addr[63924]= 1460659832;
assign addr[63925]= 1403673233;
assign addr[63926]= 1344905966;
assign addr[63927]= 1284432584;
assign addr[63928]= 1222329801;
assign addr[63929]= 1158676398;
assign addr[63930]= 1093553126;
assign addr[63931]= 1027042599;
assign addr[63932]= 959229189;
assign addr[63933]= 890198924;
assign addr[63934]= 820039373;
assign addr[63935]= 748839539;
assign addr[63936]= 676689746;
assign addr[63937]= 603681519;
assign addr[63938]= 529907477;
assign addr[63939]= 455461206;
assign addr[63940]= 380437148;
assign addr[63941]= 304930476;
assign addr[63942]= 229036977;
assign addr[63943]= 152852926;
assign addr[63944]= 76474970;
assign addr[63945]= 0;
assign addr[63946]= -76474970;
assign addr[63947]= -152852926;
assign addr[63948]= -229036977;
assign addr[63949]= -304930476;
assign addr[63950]= -380437148;
assign addr[63951]= -455461206;
assign addr[63952]= -529907477;
assign addr[63953]= -603681519;
assign addr[63954]= -676689746;
assign addr[63955]= -748839539;
assign addr[63956]= -820039373;
assign addr[63957]= -890198924;
assign addr[63958]= -959229189;
assign addr[63959]= -1027042599;
assign addr[63960]= -1093553126;
assign addr[63961]= -1158676398;
assign addr[63962]= -1222329801;
assign addr[63963]= -1284432584;
assign addr[63964]= -1344905966;
assign addr[63965]= -1403673233;
assign addr[63966]= -1460659832;
assign addr[63967]= -1515793473;
assign addr[63968]= -1569004214;
assign addr[63969]= -1620224553;
assign addr[63970]= -1669389513;
assign addr[63971]= -1716436725;
assign addr[63972]= -1761306505;
assign addr[63973]= -1803941934;
assign addr[63974]= -1844288924;
assign addr[63975]= -1882296293;
assign addr[63976]= -1917915825;
assign addr[63977]= -1951102334;
assign addr[63978]= -1981813720;
assign addr[63979]= -2010011024;
assign addr[63980]= -2035658475;
assign addr[63981]= -2058723538;
assign addr[63982]= -2079176953;
assign addr[63983]= -2096992772;
assign addr[63984]= -2112148396;
assign addr[63985]= -2124624598;
assign addr[63986]= -2134405552;
assign addr[63987]= -2141478848;
assign addr[63988]= -2145835515;
assign addr[63989]= -2147470025;
assign addr[63990]= -2146380306;
assign addr[63991]= -2142567738;
assign addr[63992]= -2136037160;
assign addr[63993]= -2126796855;
assign addr[63994]= -2114858546;
assign addr[63995]= -2100237377;
assign addr[63996]= -2082951896;
assign addr[63997]= -2063024031;
assign addr[63998]= -2040479063;
assign addr[63999]= -2015345591;
assign addr[64000]= -1987655498;
assign addr[64001]= -1957443913;
assign addr[64002]= -1924749160;
assign addr[64003]= -1889612716;
assign addr[64004]= -1852079154;
assign addr[64005]= -1812196087;
assign addr[64006]= -1770014111;
assign addr[64007]= -1725586737;
assign addr[64008]= -1678970324;
assign addr[64009]= -1630224009;
assign addr[64010]= -1579409630;
assign addr[64011]= -1526591649;
assign addr[64012]= -1471837070;
assign addr[64013]= -1415215352;
assign addr[64014]= -1356798326;
assign addr[64015]= -1296660098;
assign addr[64016]= -1234876957;
assign addr[64017]= -1171527280;
assign addr[64018]= -1106691431;
assign addr[64019]= -1040451659;
assign addr[64020]= -972891995;
assign addr[64021]= -904098143;
assign addr[64022]= -834157373;
assign addr[64023]= -763158411;
assign addr[64024]= -691191324;
assign addr[64025]= -618347408;
assign addr[64026]= -544719071;
assign addr[64027]= -470399716;
assign addr[64028]= -395483624;
assign addr[64029]= -320065829;
assign addr[64030]= -244242007;
assign addr[64031]= -168108346;
assign addr[64032]= -91761426;
assign addr[64033]= -15298099;
assign addr[64034]= 61184634;
assign addr[64035]= 137589750;
assign addr[64036]= 213820322;
assign addr[64037]= 289779648;
assign addr[64038]= 365371365;
assign addr[64039]= 440499581;
assign addr[64040]= 515068990;
assign addr[64041]= 588984994;
assign addr[64042]= 662153826;
assign addr[64043]= 734482665;
assign addr[64044]= 805879757;
assign addr[64045]= 876254528;
assign addr[64046]= 945517704;
assign addr[64047]= 1013581418;
assign addr[64048]= 1080359326;
assign addr[64049]= 1145766716;
assign addr[64050]= 1209720613;
assign addr[64051]= 1272139887;
assign addr[64052]= 1332945355;
assign addr[64053]= 1392059879;
assign addr[64054]= 1449408469;
assign addr[64055]= 1504918373;
assign addr[64056]= 1558519173;
assign addr[64057]= 1610142873;
assign addr[64058]= 1659723983;
assign addr[64059]= 1707199606;
assign addr[64060]= 1752509516;
assign addr[64061]= 1795596234;
assign addr[64062]= 1836405100;
assign addr[64063]= 1874884346;
assign addr[64064]= 1910985158;
assign addr[64065]= 1944661739;
assign addr[64066]= 1975871368;
assign addr[64067]= 2004574453;
assign addr[64068]= 2030734582;
assign addr[64069]= 2054318569;
assign addr[64070]= 2075296495;
assign addr[64071]= 2093641749;
assign addr[64072]= 2109331059;
assign addr[64073]= 2122344521;
assign addr[64074]= 2132665626;
assign addr[64075]= 2140281282;
assign addr[64076]= 2145181827;
assign addr[64077]= 2147361045;
assign addr[64078]= 2146816171;
assign addr[64079]= 2143547897;
assign addr[64080]= 2137560369;
assign addr[64081]= 2128861181;
assign addr[64082]= 2117461370;
assign addr[64083]= 2103375398;
assign addr[64084]= 2086621133;
assign addr[64085]= 2067219829;
assign addr[64086]= 2045196100;
assign addr[64087]= 2020577882;
assign addr[64088]= 1993396407;
assign addr[64089]= 1963686155;
assign addr[64090]= 1931484818;
assign addr[64091]= 1896833245;
assign addr[64092]= 1859775393;
assign addr[64093]= 1820358275;
assign addr[64094]= 1778631892;
assign addr[64095]= 1734649179;
assign addr[64096]= 1688465931;
assign addr[64097]= 1640140734;
assign addr[64098]= 1589734894;
assign addr[64099]= 1537312353;
assign addr[64100]= 1482939614;
assign addr[64101]= 1426685652;
assign addr[64102]= 1368621831;
assign addr[64103]= 1308821808;
assign addr[64104]= 1247361445;
assign addr[64105]= 1184318708;
assign addr[64106]= 1119773573;
assign addr[64107]= 1053807919;
assign addr[64108]= 986505429;
assign addr[64109]= 917951481;
assign addr[64110]= 848233042;
assign addr[64111]= 777438554;
assign addr[64112]= 705657826;
assign addr[64113]= 632981917;
assign addr[64114]= 559503022;
assign addr[64115]= 485314355;
assign addr[64116]= 410510029;
assign addr[64117]= 335184940;
assign addr[64118]= 259434643;
assign addr[64119]= 183355234;
assign addr[64120]= 107043224;
assign addr[64121]= 30595422;
assign addr[64122]= -45891193;
assign addr[64123]= -122319591;
assign addr[64124]= -198592817;
assign addr[64125]= -274614114;
assign addr[64126]= -350287041;
assign addr[64127]= -425515602;
assign addr[64128]= -500204365;
assign addr[64129]= -574258580;
assign addr[64130]= -647584304;
assign addr[64131]= -720088517;
assign addr[64132]= -791679244;
assign addr[64133]= -862265664;
assign addr[64134]= -931758235;
assign addr[64135]= -1000068799;
assign addr[64136]= -1067110699;
assign addr[64137]= -1132798888;
assign addr[64138]= -1197050035;
assign addr[64139]= -1259782632;
assign addr[64140]= -1320917099;
assign addr[64141]= -1380375881;
assign addr[64142]= -1438083551;
assign addr[64143]= -1493966902;
assign addr[64144]= -1547955041;
assign addr[64145]= -1599979481;
assign addr[64146]= -1649974225;
assign addr[64147]= -1697875851;
assign addr[64148]= -1743623590;
assign addr[64149]= -1787159411;
assign addr[64150]= -1828428082;
assign addr[64151]= -1867377253;
assign addr[64152]= -1903957513;
assign addr[64153]= -1938122457;
assign addr[64154]= -1969828744;
assign addr[64155]= -1999036154;
assign addr[64156]= -2025707632;
assign addr[64157]= -2049809346;
assign addr[64158]= -2071310720;
assign addr[64159]= -2090184478;
assign addr[64160]= -2106406677;
assign addr[64161]= -2119956737;
assign addr[64162]= -2130817471;
assign addr[64163]= -2138975100;
assign addr[64164]= -2144419275;
assign addr[64165]= -2147143090;
assign addr[64166]= -2147143090;
assign addr[64167]= -2144419275;
assign addr[64168]= -2138975100;
assign addr[64169]= -2130817471;
assign addr[64170]= -2119956737;
assign addr[64171]= -2106406677;
assign addr[64172]= -2090184478;
assign addr[64173]= -2071310720;
assign addr[64174]= -2049809346;
assign addr[64175]= -2025707632;
assign addr[64176]= -1999036154;
assign addr[64177]= -1969828744;
assign addr[64178]= -1938122457;
assign addr[64179]= -1903957513;
assign addr[64180]= -1867377253;
assign addr[64181]= -1828428082;
assign addr[64182]= -1787159411;
assign addr[64183]= -1743623590;
assign addr[64184]= -1697875851;
assign addr[64185]= -1649974225;
assign addr[64186]= -1599979481;
assign addr[64187]= -1547955041;
assign addr[64188]= -1493966902;
assign addr[64189]= -1438083551;
assign addr[64190]= -1380375881;
assign addr[64191]= -1320917099;
assign addr[64192]= -1259782632;
assign addr[64193]= -1197050035;
assign addr[64194]= -1132798888;
assign addr[64195]= -1067110699;
assign addr[64196]= -1000068799;
assign addr[64197]= -931758235;
assign addr[64198]= -862265664;
assign addr[64199]= -791679244;
assign addr[64200]= -720088517;
assign addr[64201]= -647584304;
assign addr[64202]= -574258580;
assign addr[64203]= -500204365;
assign addr[64204]= -425515602;
assign addr[64205]= -350287041;
assign addr[64206]= -274614114;
assign addr[64207]= -198592817;
assign addr[64208]= -122319591;
assign addr[64209]= -45891193;
assign addr[64210]= 30595422;
assign addr[64211]= 107043224;
assign addr[64212]= 183355234;
assign addr[64213]= 259434643;
assign addr[64214]= 335184940;
assign addr[64215]= 410510029;
assign addr[64216]= 485314355;
assign addr[64217]= 559503022;
assign addr[64218]= 632981917;
assign addr[64219]= 705657826;
assign addr[64220]= 777438554;
assign addr[64221]= 848233042;
assign addr[64222]= 917951481;
assign addr[64223]= 986505429;
assign addr[64224]= 1053807919;
assign addr[64225]= 1119773573;
assign addr[64226]= 1184318708;
assign addr[64227]= 1247361445;
assign addr[64228]= 1308821808;
assign addr[64229]= 1368621831;
assign addr[64230]= 1426685652;
assign addr[64231]= 1482939614;
assign addr[64232]= 1537312353;
assign addr[64233]= 1589734894;
assign addr[64234]= 1640140734;
assign addr[64235]= 1688465931;
assign addr[64236]= 1734649179;
assign addr[64237]= 1778631892;
assign addr[64238]= 1820358275;
assign addr[64239]= 1859775393;
assign addr[64240]= 1896833245;
assign addr[64241]= 1931484818;
assign addr[64242]= 1963686155;
assign addr[64243]= 1993396407;
assign addr[64244]= 2020577882;
assign addr[64245]= 2045196100;
assign addr[64246]= 2067219829;
assign addr[64247]= 2086621133;
assign addr[64248]= 2103375398;
assign addr[64249]= 2117461370;
assign addr[64250]= 2128861181;
assign addr[64251]= 2137560369;
assign addr[64252]= 2143547897;
assign addr[64253]= 2146816171;
assign addr[64254]= 2147361045;
assign addr[64255]= 2145181827;
assign addr[64256]= 2140281282;
assign addr[64257]= 2132665626;
assign addr[64258]= 2122344521;
assign addr[64259]= 2109331059;
assign addr[64260]= 2093641749;
assign addr[64261]= 2075296495;
assign addr[64262]= 2054318569;
assign addr[64263]= 2030734582;
assign addr[64264]= 2004574453;
assign addr[64265]= 1975871368;
assign addr[64266]= 1944661739;
assign addr[64267]= 1910985158;
assign addr[64268]= 1874884346;
assign addr[64269]= 1836405100;
assign addr[64270]= 1795596234;
assign addr[64271]= 1752509516;
assign addr[64272]= 1707199606;
assign addr[64273]= 1659723983;
assign addr[64274]= 1610142873;
assign addr[64275]= 1558519173;
assign addr[64276]= 1504918373;
assign addr[64277]= 1449408469;
assign addr[64278]= 1392059879;
assign addr[64279]= 1332945355;
assign addr[64280]= 1272139887;
assign addr[64281]= 1209720613;
assign addr[64282]= 1145766716;
assign addr[64283]= 1080359326;
assign addr[64284]= 1013581418;
assign addr[64285]= 945517704;
assign addr[64286]= 876254528;
assign addr[64287]= 805879757;
assign addr[64288]= 734482665;
assign addr[64289]= 662153826;
assign addr[64290]= 588984994;
assign addr[64291]= 515068990;
assign addr[64292]= 440499581;
assign addr[64293]= 365371365;
assign addr[64294]= 289779648;
assign addr[64295]= 213820322;
assign addr[64296]= 137589750;
assign addr[64297]= 61184634;
assign addr[64298]= -15298099;
assign addr[64299]= -91761426;
assign addr[64300]= -168108346;
assign addr[64301]= -244242007;
assign addr[64302]= -320065829;
assign addr[64303]= -395483624;
assign addr[64304]= -470399716;
assign addr[64305]= -544719071;
assign addr[64306]= -618347408;
assign addr[64307]= -691191324;
assign addr[64308]= -763158411;
assign addr[64309]= -834157373;
assign addr[64310]= -904098143;
assign addr[64311]= -972891995;
assign addr[64312]= -1040451659;
assign addr[64313]= -1106691431;
assign addr[64314]= -1171527280;
assign addr[64315]= -1234876957;
assign addr[64316]= -1296660098;
assign addr[64317]= -1356798326;
assign addr[64318]= -1415215352;
assign addr[64319]= -1471837070;
assign addr[64320]= -1526591649;
assign addr[64321]= -1579409630;
assign addr[64322]= -1630224009;
assign addr[64323]= -1678970324;
assign addr[64324]= -1725586737;
assign addr[64325]= -1770014111;
assign addr[64326]= -1812196087;
assign addr[64327]= -1852079154;
assign addr[64328]= -1889612716;
assign addr[64329]= -1924749160;
assign addr[64330]= -1957443913;
assign addr[64331]= -1987655498;
assign addr[64332]= -2015345591;
assign addr[64333]= -2040479063;
assign addr[64334]= -2063024031;
assign addr[64335]= -2082951896;
assign addr[64336]= -2100237377;
assign addr[64337]= -2114858546;
assign addr[64338]= -2126796855;
assign addr[64339]= -2136037160;
assign addr[64340]= -2142567738;
assign addr[64341]= -2146380306;
assign addr[64342]= -2147470025;
assign addr[64343]= -2145835515;
assign addr[64344]= -2141478848;
assign addr[64345]= -2134405552;
assign addr[64346]= -2124624598;
assign addr[64347]= -2112148396;
assign addr[64348]= -2096992772;
assign addr[64349]= -2079176953;
assign addr[64350]= -2058723538;
assign addr[64351]= -2035658475;
assign addr[64352]= -2010011024;
assign addr[64353]= -1981813720;
assign addr[64354]= -1951102334;
assign addr[64355]= -1917915825;
assign addr[64356]= -1882296293;
assign addr[64357]= -1844288924;
assign addr[64358]= -1803941934;
assign addr[64359]= -1761306505;
assign addr[64360]= -1716436725;
assign addr[64361]= -1669389513;
assign addr[64362]= -1620224553;
assign addr[64363]= -1569004214;
assign addr[64364]= -1515793473;
assign addr[64365]= -1460659832;
assign addr[64366]= -1403673233;
assign addr[64367]= -1344905966;
assign addr[64368]= -1284432584;
assign addr[64369]= -1222329801;
assign addr[64370]= -1158676398;
assign addr[64371]= -1093553126;
assign addr[64372]= -1027042599;
assign addr[64373]= -959229189;
assign addr[64374]= -890198924;
assign addr[64375]= -820039373;
assign addr[64376]= -748839539;
assign addr[64377]= -676689746;
assign addr[64378]= -603681519;
assign addr[64379]= -529907477;
assign addr[64380]= -455461206;
assign addr[64381]= -380437148;
assign addr[64382]= -304930476;
assign addr[64383]= -229036977;
assign addr[64384]= -152852926;
assign addr[64385]= -76474970;
assign addr[64386]= 0;
assign addr[64387]= 76474970;
assign addr[64388]= 152852926;
assign addr[64389]= 229036977;
assign addr[64390]= 304930476;
assign addr[64391]= 380437148;
assign addr[64392]= 455461206;
assign addr[64393]= 529907477;
assign addr[64394]= 603681519;
assign addr[64395]= 676689746;
assign addr[64396]= 748839539;
assign addr[64397]= 820039373;
assign addr[64398]= 890198924;
assign addr[64399]= 959229189;
assign addr[64400]= 1027042599;
assign addr[64401]= 1093553126;
assign addr[64402]= 1158676398;
assign addr[64403]= 1222329801;
assign addr[64404]= 1284432584;
assign addr[64405]= 1344905966;
assign addr[64406]= 1403673233;
assign addr[64407]= 1460659832;
assign addr[64408]= 1515793473;
assign addr[64409]= 1569004214;
assign addr[64410]= 1620224553;
assign addr[64411]= 1669389513;
assign addr[64412]= 1716436725;
assign addr[64413]= 1761306505;
assign addr[64414]= 1803941934;
assign addr[64415]= 1844288924;
assign addr[64416]= 1882296293;
assign addr[64417]= 1917915825;
assign addr[64418]= 1951102334;
assign addr[64419]= 1981813720;
assign addr[64420]= 2010011024;
assign addr[64421]= 2035658475;
assign addr[64422]= 2058723538;
assign addr[64423]= 2079176953;
assign addr[64424]= 2096992772;
assign addr[64425]= 2112148396;
assign addr[64426]= 2124624598;
assign addr[64427]= 2134405552;
assign addr[64428]= 2141478848;
assign addr[64429]= 2145835515;
assign addr[64430]= 2147470025;
assign addr[64431]= 2146380306;
assign addr[64432]= 2142567738;
assign addr[64433]= 2136037160;
assign addr[64434]= 2126796855;
assign addr[64435]= 2114858546;
assign addr[64436]= 2100237377;
assign addr[64437]= 2082951896;
assign addr[64438]= 2063024031;
assign addr[64439]= 2040479063;
assign addr[64440]= 2015345591;
assign addr[64441]= 1987655498;
assign addr[64442]= 1957443913;
assign addr[64443]= 1924749160;
assign addr[64444]= 1889612716;
assign addr[64445]= 1852079154;
assign addr[64446]= 1812196087;
assign addr[64447]= 1770014111;
assign addr[64448]= 1725586737;
assign addr[64449]= 1678970324;
assign addr[64450]= 1630224009;
assign addr[64451]= 1579409630;
assign addr[64452]= 1526591649;
assign addr[64453]= 1471837070;
assign addr[64454]= 1415215352;
assign addr[64455]= 1356798326;
assign addr[64456]= 1296660098;
assign addr[64457]= 1234876957;
assign addr[64458]= 1171527280;
assign addr[64459]= 1106691431;
assign addr[64460]= 1040451659;
assign addr[64461]= 972891995;
assign addr[64462]= 904098143;
assign addr[64463]= 834157373;
assign addr[64464]= 763158411;
assign addr[64465]= 691191324;
assign addr[64466]= 618347408;
assign addr[64467]= 544719071;
assign addr[64468]= 470399716;
assign addr[64469]= 395483624;
assign addr[64470]= 320065829;
assign addr[64471]= 244242007;
assign addr[64472]= 168108346;
assign addr[64473]= 91761426;
assign addr[64474]= 15298099;
assign addr[64475]= -61184634;
assign addr[64476]= -137589750;
assign addr[64477]= -213820322;
assign addr[64478]= -289779648;
assign addr[64479]= -365371365;
assign addr[64480]= -440499581;
assign addr[64481]= -515068990;
assign addr[64482]= -588984994;
assign addr[64483]= -662153826;
assign addr[64484]= -734482665;
assign addr[64485]= -805879757;
assign addr[64486]= -876254528;
assign addr[64487]= -945517704;
assign addr[64488]= -1013581418;
assign addr[64489]= -1080359326;
assign addr[64490]= -1145766716;
assign addr[64491]= -1209720613;
assign addr[64492]= -1272139887;
assign addr[64493]= -1332945355;
assign addr[64494]= -1392059879;
assign addr[64495]= -1449408469;
assign addr[64496]= -1504918373;
assign addr[64497]= -1558519173;
assign addr[64498]= -1610142873;
assign addr[64499]= -1659723983;
assign addr[64500]= -1707199606;
assign addr[64501]= -1752509516;
assign addr[64502]= -1795596234;
assign addr[64503]= -1836405100;
assign addr[64504]= -1874884346;
assign addr[64505]= -1910985158;
assign addr[64506]= -1944661739;
assign addr[64507]= -1975871368;
assign addr[64508]= -2004574453;
assign addr[64509]= -2030734582;
assign addr[64510]= -2054318569;
assign addr[64511]= -2075296495;
assign addr[64512]= -2093641749;
assign addr[64513]= -2109331059;
assign addr[64514]= -2122344521;
assign addr[64515]= -2132665626;
assign addr[64516]= -2140281282;
assign addr[64517]= -2145181827;
assign addr[64518]= -2147361045;
assign addr[64519]= -2146816171;
assign addr[64520]= -2143547897;
assign addr[64521]= -2137560369;
assign addr[64522]= -2128861181;
assign addr[64523]= -2117461370;
assign addr[64524]= -2103375398;
assign addr[64525]= -2086621133;
assign addr[64526]= -2067219829;
assign addr[64527]= -2045196100;
assign addr[64528]= -2020577882;
assign addr[64529]= -1993396407;
assign addr[64530]= -1963686155;
assign addr[64531]= -1931484818;
assign addr[64532]= -1896833245;
assign addr[64533]= -1859775393;
assign addr[64534]= -1820358275;
assign addr[64535]= -1778631892;
assign addr[64536]= -1734649179;
assign addr[64537]= -1688465931;
assign addr[64538]= -1640140734;
assign addr[64539]= -1589734894;
assign addr[64540]= -1537312353;
assign addr[64541]= -1482939614;
assign addr[64542]= -1426685652;
assign addr[64543]= -1368621831;
assign addr[64544]= -1308821808;
assign addr[64545]= -1247361445;
assign addr[64546]= -1184318708;
assign addr[64547]= -1119773573;
assign addr[64548]= -1053807919;
assign addr[64549]= -986505429;
assign addr[64550]= -917951481;
assign addr[64551]= -848233042;
assign addr[64552]= -777438554;
assign addr[64553]= -705657826;
assign addr[64554]= -632981917;
assign addr[64555]= -559503022;
assign addr[64556]= -485314355;
assign addr[64557]= -410510029;
assign addr[64558]= -335184940;
assign addr[64559]= -259434643;
assign addr[64560]= -183355234;
assign addr[64561]= -107043224;
assign addr[64562]= -30595422;
assign addr[64563]= 45891193;
assign addr[64564]= 122319591;
assign addr[64565]= 198592817;
assign addr[64566]= 274614114;
assign addr[64567]= 350287041;
assign addr[64568]= 425515602;
assign addr[64569]= 500204365;
assign addr[64570]= 574258580;
assign addr[64571]= 647584304;
assign addr[64572]= 720088517;
assign addr[64573]= 791679244;
assign addr[64574]= 862265664;
assign addr[64575]= 931758235;
assign addr[64576]= 1000068799;
assign addr[64577]= 1067110699;
assign addr[64578]= 1132798888;
assign addr[64579]= 1197050035;
assign addr[64580]= 1259782632;
assign addr[64581]= 1320917099;
assign addr[64582]= 1380375881;
assign addr[64583]= 1438083551;
assign addr[64584]= 1493966902;
assign addr[64585]= 1547955041;
assign addr[64586]= 1599979481;
assign addr[64587]= 1649974225;
assign addr[64588]= 1697875851;
assign addr[64589]= 1743623590;
assign addr[64590]= 1787159411;
assign addr[64591]= 1828428082;
assign addr[64592]= 1867377253;
assign addr[64593]= 1903957513;
assign addr[64594]= 1938122457;
assign addr[64595]= 1969828744;
assign addr[64596]= 1999036154;
assign addr[64597]= 2025707632;
assign addr[64598]= 2049809346;
assign addr[64599]= 2071310720;
assign addr[64600]= 2090184478;
assign addr[64601]= 2106406677;
assign addr[64602]= 2119956737;
assign addr[64603]= 2130817471;
assign addr[64604]= 2138975100;
assign addr[64605]= 2144419275;
assign addr[64606]= 2147143090;
assign addr[64607]= 2147143090;
assign addr[64608]= 2144419275;
assign addr[64609]= 2138975100;
assign addr[64610]= 2130817471;
assign addr[64611]= 2119956737;
assign addr[64612]= 2106406677;
assign addr[64613]= 2090184478;
assign addr[64614]= 2071310720;
assign addr[64615]= 2049809346;
assign addr[64616]= 2025707632;
assign addr[64617]= 1999036154;
assign addr[64618]= 1969828744;
assign addr[64619]= 1938122457;
assign addr[64620]= 1903957513;
assign addr[64621]= 1867377253;
assign addr[64622]= 1828428082;
assign addr[64623]= 1787159411;
assign addr[64624]= 1743623590;
assign addr[64625]= 1697875851;
assign addr[64626]= 1649974225;
assign addr[64627]= 1599979481;
assign addr[64628]= 1547955041;
assign addr[64629]= 1493966902;
assign addr[64630]= 1438083551;
assign addr[64631]= 1380375881;
assign addr[64632]= 1320917099;
assign addr[64633]= 1259782632;
assign addr[64634]= 1197050035;
assign addr[64635]= 1132798888;
assign addr[64636]= 1067110699;
assign addr[64637]= 1000068799;
assign addr[64638]= 931758235;
assign addr[64639]= 862265664;
assign addr[64640]= 791679244;
assign addr[64641]= 720088517;
assign addr[64642]= 647584304;
assign addr[64643]= 574258580;
assign addr[64644]= 500204365;
assign addr[64645]= 425515602;
assign addr[64646]= 350287041;
assign addr[64647]= 274614114;
assign addr[64648]= 198592817;
assign addr[64649]= 122319591;
assign addr[64650]= 45891193;
assign addr[64651]= -30595422;
assign addr[64652]= -107043224;
assign addr[64653]= -183355234;
assign addr[64654]= -259434643;
assign addr[64655]= -335184940;
assign addr[64656]= -410510029;
assign addr[64657]= -485314355;
assign addr[64658]= -559503022;
assign addr[64659]= -632981917;
assign addr[64660]= -705657826;
assign addr[64661]= -777438554;
assign addr[64662]= -848233042;
assign addr[64663]= -917951481;
assign addr[64664]= -986505429;
assign addr[64665]= -1053807919;
assign addr[64666]= -1119773573;
assign addr[64667]= -1184318708;
assign addr[64668]= -1247361445;
assign addr[64669]= -1308821808;
assign addr[64670]= -1368621831;
assign addr[64671]= -1426685652;
assign addr[64672]= -1482939614;
assign addr[64673]= -1537312353;
assign addr[64674]= -1589734894;
assign addr[64675]= -1640140734;
assign addr[64676]= -1688465931;
assign addr[64677]= -1734649179;
assign addr[64678]= -1778631892;
assign addr[64679]= -1820358275;
assign addr[64680]= -1859775393;
assign addr[64681]= -1896833245;
assign addr[64682]= -1931484818;
assign addr[64683]= -1963686155;
assign addr[64684]= -1993396407;
assign addr[64685]= -2020577882;
assign addr[64686]= -2045196100;
assign addr[64687]= -2067219829;
assign addr[64688]= -2086621133;
assign addr[64689]= -2103375398;
assign addr[64690]= -2117461370;
assign addr[64691]= -2128861181;
assign addr[64692]= -2137560369;
assign addr[64693]= -2143547897;
assign addr[64694]= -2146816171;
assign addr[64695]= -2147361045;
assign addr[64696]= -2145181827;
assign addr[64697]= -2140281282;
assign addr[64698]= -2132665626;
assign addr[64699]= -2122344521;
assign addr[64700]= -2109331059;
assign addr[64701]= -2093641749;
assign addr[64702]= -2075296495;
assign addr[64703]= -2054318569;
assign addr[64704]= -2030734582;
assign addr[64705]= -2004574453;
assign addr[64706]= -1975871368;
assign addr[64707]= -1944661739;
assign addr[64708]= -1910985158;
assign addr[64709]= -1874884346;
assign addr[64710]= -1836405100;
assign addr[64711]= -1795596234;
assign addr[64712]= -1752509516;
assign addr[64713]= -1707199606;
assign addr[64714]= -1659723983;
assign addr[64715]= -1610142873;
assign addr[64716]= -1558519173;
assign addr[64717]= -1504918373;
assign addr[64718]= -1449408469;
assign addr[64719]= -1392059879;
assign addr[64720]= -1332945355;
assign addr[64721]= -1272139887;
assign addr[64722]= -1209720613;
assign addr[64723]= -1145766716;
assign addr[64724]= -1080359326;
assign addr[64725]= -1013581418;
assign addr[64726]= -945517704;
assign addr[64727]= -876254528;
assign addr[64728]= -805879757;
assign addr[64729]= -734482665;
assign addr[64730]= -662153826;
assign addr[64731]= -588984994;
assign addr[64732]= -515068990;
assign addr[64733]= -440499581;
assign addr[64734]= -365371365;
assign addr[64735]= -289779648;
assign addr[64736]= -213820322;
assign addr[64737]= -137589750;
assign addr[64738]= -61184634;
assign addr[64739]= 15298099;
assign addr[64740]= 91761426;
assign addr[64741]= 168108346;
assign addr[64742]= 244242007;
assign addr[64743]= 320065829;
assign addr[64744]= 395483624;
assign addr[64745]= 470399716;
assign addr[64746]= 544719071;
assign addr[64747]= 618347408;
assign addr[64748]= 691191324;
assign addr[64749]= 763158411;
assign addr[64750]= 834157373;
assign addr[64751]= 904098143;
assign addr[64752]= 972891995;
assign addr[64753]= 1040451659;
assign addr[64754]= 1106691431;
assign addr[64755]= 1171527280;
assign addr[64756]= 1234876957;
assign addr[64757]= 1296660098;
assign addr[64758]= 1356798326;
assign addr[64759]= 1415215352;
assign addr[64760]= 1471837070;
assign addr[64761]= 1526591649;
assign addr[64762]= 1579409630;
assign addr[64763]= 1630224009;
assign addr[64764]= 1678970324;
assign addr[64765]= 1725586737;
assign addr[64766]= 1770014111;
assign addr[64767]= 1812196087;
assign addr[64768]= 1852079154;
assign addr[64769]= 1889612716;
assign addr[64770]= 1924749160;
assign addr[64771]= 1957443913;
assign addr[64772]= 1987655498;
assign addr[64773]= 2015345591;
assign addr[64774]= 2040479063;
assign addr[64775]= 2063024031;
assign addr[64776]= 2082951896;
assign addr[64777]= 2100237377;
assign addr[64778]= 2114858546;
assign addr[64779]= 2126796855;
assign addr[64780]= 2136037160;
assign addr[64781]= 2142567738;
assign addr[64782]= 2146380306;
assign addr[64783]= 2147470025;
assign addr[64784]= 2145835515;
assign addr[64785]= 2141478848;
assign addr[64786]= 2134405552;
assign addr[64787]= 2124624598;
assign addr[64788]= 2112148396;
assign addr[64789]= 2096992772;
assign addr[64790]= 2079176953;
assign addr[64791]= 2058723538;
assign addr[64792]= 2035658475;
assign addr[64793]= 2010011024;
assign addr[64794]= 1981813720;
assign addr[64795]= 1951102334;
assign addr[64796]= 1917915825;
assign addr[64797]= 1882296293;
assign addr[64798]= 1844288924;
assign addr[64799]= 1803941934;
assign addr[64800]= 1761306505;
assign addr[64801]= 1716436725;
assign addr[64802]= 1669389513;
assign addr[64803]= 1620224553;
assign addr[64804]= 1569004214;
assign addr[64805]= 1515793473;
assign addr[64806]= 1460659832;
assign addr[64807]= 1403673233;
assign addr[64808]= 1344905966;
assign addr[64809]= 1284432584;
assign addr[64810]= 1222329801;
assign addr[64811]= 1158676398;
assign addr[64812]= 1093553126;
assign addr[64813]= 1027042599;
assign addr[64814]= 959229189;
assign addr[64815]= 890198924;
assign addr[64816]= 820039373;
assign addr[64817]= 748839539;
assign addr[64818]= 676689746;
assign addr[64819]= 603681519;
assign addr[64820]= 529907477;
assign addr[64821]= 455461206;
assign addr[64822]= 380437148;
assign addr[64823]= 304930476;
assign addr[64824]= 229036977;
assign addr[64825]= 152852926;
assign addr[64826]= 76474970;
assign addr[64827]= 0;
assign addr[64828]= -76474970;
assign addr[64829]= -152852926;
assign addr[64830]= -229036977;
assign addr[64831]= -304930476;
assign addr[64832]= -380437148;
assign addr[64833]= -455461206;
assign addr[64834]= -529907477;
assign addr[64835]= -603681519;
assign addr[64836]= -676689746;
assign addr[64837]= -748839539;
assign addr[64838]= -820039373;
assign addr[64839]= -890198924;
assign addr[64840]= -959229189;
assign addr[64841]= -1027042599;
assign addr[64842]= -1093553126;
assign addr[64843]= -1158676398;
assign addr[64844]= -1222329801;
assign addr[64845]= -1284432584;
assign addr[64846]= -1344905966;
assign addr[64847]= -1403673233;
assign addr[64848]= -1460659832;
assign addr[64849]= -1515793473;
assign addr[64850]= -1569004214;
assign addr[64851]= -1620224553;
assign addr[64852]= -1669389513;
assign addr[64853]= -1716436725;
assign addr[64854]= -1761306505;
assign addr[64855]= -1803941934;
assign addr[64856]= -1844288924;
assign addr[64857]= -1882296293;
assign addr[64858]= -1917915825;
assign addr[64859]= -1951102334;
assign addr[64860]= -1981813720;
assign addr[64861]= -2010011024;
assign addr[64862]= -2035658475;
assign addr[64863]= -2058723538;
assign addr[64864]= -2079176953;
assign addr[64865]= -2096992772;
assign addr[64866]= -2112148396;
assign addr[64867]= -2124624598;
assign addr[64868]= -2134405552;
assign addr[64869]= -2141478848;
assign addr[64870]= -2145835515;
assign addr[64871]= -2147470025;
assign addr[64872]= -2146380306;
assign addr[64873]= -2142567738;
assign addr[64874]= -2136037160;
assign addr[64875]= -2126796855;
assign addr[64876]= -2114858546;
assign addr[64877]= -2100237377;
assign addr[64878]= -2082951896;
assign addr[64879]= -2063024031;
assign addr[64880]= -2040479063;
assign addr[64881]= -2015345591;
assign addr[64882]= -1987655498;
assign addr[64883]= -1957443913;
assign addr[64884]= -1924749160;
assign addr[64885]= -1889612716;
assign addr[64886]= -1852079154;
assign addr[64887]= -1812196087;
assign addr[64888]= -1770014111;
assign addr[64889]= -1725586737;
assign addr[64890]= -1678970324;
assign addr[64891]= -1630224009;
assign addr[64892]= -1579409630;
assign addr[64893]= -1526591649;
assign addr[64894]= -1471837070;
assign addr[64895]= -1415215352;
assign addr[64896]= -1356798326;
assign addr[64897]= -1296660098;
assign addr[64898]= -1234876957;
assign addr[64899]= -1171527280;
assign addr[64900]= -1106691431;
assign addr[64901]= -1040451659;
assign addr[64902]= -972891995;
assign addr[64903]= -904098143;
assign addr[64904]= -834157373;
assign addr[64905]= -763158411;
assign addr[64906]= -691191324;
assign addr[64907]= -618347408;
assign addr[64908]= -544719071;
assign addr[64909]= -470399716;
assign addr[64910]= -395483624;
assign addr[64911]= -320065829;
assign addr[64912]= -244242007;
assign addr[64913]= -168108346;
assign addr[64914]= -91761426;
assign addr[64915]= -15298099;
assign addr[64916]= 61184634;
assign addr[64917]= 137589750;
assign addr[64918]= 213820322;
assign addr[64919]= 289779648;
assign addr[64920]= 365371365;
assign addr[64921]= 440499581;
assign addr[64922]= 515068990;
assign addr[64923]= 588984994;
assign addr[64924]= 662153826;
assign addr[64925]= 734482665;
assign addr[64926]= 805879757;
assign addr[64927]= 876254528;
assign addr[64928]= 945517704;
assign addr[64929]= 1013581418;
assign addr[64930]= 1080359326;
assign addr[64931]= 1145766716;
assign addr[64932]= 1209720613;
assign addr[64933]= 1272139887;
assign addr[64934]= 1332945355;
assign addr[64935]= 1392059879;
assign addr[64936]= 1449408469;
assign addr[64937]= 1504918373;
assign addr[64938]= 1558519173;
assign addr[64939]= 1610142873;
assign addr[64940]= 1659723983;
assign addr[64941]= 1707199606;
assign addr[64942]= 1752509516;
assign addr[64943]= 1795596234;
assign addr[64944]= 1836405100;
assign addr[64945]= 1874884346;
assign addr[64946]= 1910985158;
assign addr[64947]= 1944661739;
assign addr[64948]= 1975871368;
assign addr[64949]= 2004574453;
assign addr[64950]= 2030734582;
assign addr[64951]= 2054318569;
assign addr[64952]= 2075296495;
assign addr[64953]= 2093641749;
assign addr[64954]= 2109331059;
assign addr[64955]= 2122344521;
assign addr[64956]= 2132665626;
assign addr[64957]= 2140281282;
assign addr[64958]= 2145181827;
assign addr[64959]= 2147361045;
assign addr[64960]= 2146816171;
assign addr[64961]= 2143547897;
assign addr[64962]= 2137560369;
assign addr[64963]= 2128861181;
assign addr[64964]= 2117461370;
assign addr[64965]= 2103375398;
assign addr[64966]= 2086621133;
assign addr[64967]= 2067219829;
assign addr[64968]= 2045196100;
assign addr[64969]= 2020577882;
assign addr[64970]= 1993396407;
assign addr[64971]= 1963686155;
assign addr[64972]= 1931484818;
assign addr[64973]= 1896833245;
assign addr[64974]= 1859775393;
assign addr[64975]= 1820358275;
assign addr[64976]= 1778631892;
assign addr[64977]= 1734649179;
assign addr[64978]= 1688465931;
assign addr[64979]= 1640140734;
assign addr[64980]= 1589734894;
assign addr[64981]= 1537312353;
assign addr[64982]= 1482939614;
assign addr[64983]= 1426685652;
assign addr[64984]= 1368621831;
assign addr[64985]= 1308821808;
assign addr[64986]= 1247361445;
assign addr[64987]= 1184318708;
assign addr[64988]= 1119773573;
assign addr[64989]= 1053807919;
assign addr[64990]= 986505429;
assign addr[64991]= 917951481;
assign addr[64992]= 848233042;
assign addr[64993]= 777438554;
assign addr[64994]= 705657826;
assign addr[64995]= 632981917;
assign addr[64996]= 559503022;
assign addr[64997]= 485314355;
assign addr[64998]= 410510029;
assign addr[64999]= 335184940;
assign addr[65000]= 259434643;
assign addr[65001]= 183355234;
assign addr[65002]= 107043224;
assign addr[65003]= 30595422;
assign addr[65004]= -45891193;
assign addr[65005]= -122319591;
assign addr[65006]= -198592817;
assign addr[65007]= -274614114;
assign addr[65008]= -350287041;
assign addr[65009]= -425515602;
assign addr[65010]= -500204365;
assign addr[65011]= -574258580;
assign addr[65012]= -647584304;
assign addr[65013]= -720088517;
assign addr[65014]= -791679244;
assign addr[65015]= -862265664;
assign addr[65016]= -931758235;
assign addr[65017]= -1000068799;
assign addr[65018]= -1067110699;
assign addr[65019]= -1132798888;
assign addr[65020]= -1197050035;
assign addr[65021]= -1259782632;
assign addr[65022]= -1320917099;
assign addr[65023]= -1380375881;
assign addr[65024]= -1438083551;
assign addr[65025]= -1493966902;
assign addr[65026]= -1547955041;
assign addr[65027]= -1599979481;
assign addr[65028]= -1649974225;
assign addr[65029]= -1697875851;
assign addr[65030]= -1743623590;
assign addr[65031]= -1787159411;
assign addr[65032]= -1828428082;
assign addr[65033]= -1867377253;
assign addr[65034]= -1903957513;
assign addr[65035]= -1938122457;
assign addr[65036]= -1969828744;
assign addr[65037]= -1999036154;
assign addr[65038]= -2025707632;
assign addr[65039]= -2049809346;
assign addr[65040]= -2071310720;
assign addr[65041]= -2090184478;
assign addr[65042]= -2106406677;
assign addr[65043]= -2119956737;
assign addr[65044]= -2130817471;
assign addr[65045]= -2138975100;
assign addr[65046]= -2144419275;
assign addr[65047]= -2147143090;
assign addr[65048]= -2147143090;
assign addr[65049]= -2144419275;
assign addr[65050]= -2138975100;
assign addr[65051]= -2130817471;
assign addr[65052]= -2119956737;
assign addr[65053]= -2106406677;
assign addr[65054]= -2090184478;
assign addr[65055]= -2071310720;
assign addr[65056]= -2049809346;
assign addr[65057]= -2025707632;
assign addr[65058]= -1999036154;
assign addr[65059]= -1969828744;
assign addr[65060]= -1938122457;
assign addr[65061]= -1903957513;
assign addr[65062]= -1867377253;
assign addr[65063]= -1828428082;
assign addr[65064]= -1787159411;
assign addr[65065]= -1743623590;
assign addr[65066]= -1697875851;
assign addr[65067]= -1649974225;
assign addr[65068]= -1599979481;
assign addr[65069]= -1547955041;
assign addr[65070]= -1493966902;
assign addr[65071]= -1438083551;
assign addr[65072]= -1380375881;
assign addr[65073]= -1320917099;
assign addr[65074]= -1259782632;
assign addr[65075]= -1197050035;
assign addr[65076]= -1132798888;
assign addr[65077]= -1067110699;
assign addr[65078]= -1000068799;
assign addr[65079]= -931758235;
assign addr[65080]= -862265664;
assign addr[65081]= -791679244;
assign addr[65082]= -720088517;
assign addr[65083]= -647584304;
assign addr[65084]= -574258580;
assign addr[65085]= -500204365;
assign addr[65086]= -425515602;
assign addr[65087]= -350287041;
assign addr[65088]= -274614114;
assign addr[65089]= -198592817;
assign addr[65090]= -122319591;
assign addr[65091]= -45891193;
assign addr[65092]= 30595422;
assign addr[65093]= 107043224;
assign addr[65094]= 183355234;
assign addr[65095]= 259434643;
assign addr[65096]= 335184940;
assign addr[65097]= 410510029;
assign addr[65098]= 485314355;
assign addr[65099]= 559503022;
assign addr[65100]= 632981917;
assign addr[65101]= 705657826;
assign addr[65102]= 777438554;
assign addr[65103]= 848233042;
assign addr[65104]= 917951481;
assign addr[65105]= 986505429;
assign addr[65106]= 1053807919;
assign addr[65107]= 1119773573;
assign addr[65108]= 1184318708;
assign addr[65109]= 1247361445;
assign addr[65110]= 1308821808;
assign addr[65111]= 1368621831;
assign addr[65112]= 1426685652;
assign addr[65113]= 1482939614;
assign addr[65114]= 1537312353;
assign addr[65115]= 1589734894;
assign addr[65116]= 1640140734;
assign addr[65117]= 1688465931;
assign addr[65118]= 1734649179;
assign addr[65119]= 1778631892;
assign addr[65120]= 1820358275;
assign addr[65121]= 1859775393;
assign addr[65122]= 1896833245;
assign addr[65123]= 1931484818;
assign addr[65124]= 1963686155;
assign addr[65125]= 1993396407;
assign addr[65126]= 2020577882;
assign addr[65127]= 2045196100;
assign addr[65128]= 2067219829;
assign addr[65129]= 2086621133;
assign addr[65130]= 2103375398;
assign addr[65131]= 2117461370;
assign addr[65132]= 2128861181;
assign addr[65133]= 2137560369;
assign addr[65134]= 2143547897;
assign addr[65135]= 2146816171;
assign addr[65136]= 2147361045;
assign addr[65137]= 2145181827;
assign addr[65138]= 2140281282;
assign addr[65139]= 2132665626;
assign addr[65140]= 2122344521;
assign addr[65141]= 2109331059;
assign addr[65142]= 2093641749;
assign addr[65143]= 2075296495;
assign addr[65144]= 2054318569;
assign addr[65145]= 2030734582;
assign addr[65146]= 2004574453;
assign addr[65147]= 1975871368;
assign addr[65148]= 1944661739;
assign addr[65149]= 1910985158;
assign addr[65150]= 1874884346;
assign addr[65151]= 1836405100;
assign addr[65152]= 1795596234;
assign addr[65153]= 1752509516;
assign addr[65154]= 1707199606;
assign addr[65155]= 1659723983;
assign addr[65156]= 1610142873;
assign addr[65157]= 1558519173;
assign addr[65158]= 1504918373;
assign addr[65159]= 1449408469;
assign addr[65160]= 1392059879;
assign addr[65161]= 1332945355;
assign addr[65162]= 1272139887;
assign addr[65163]= 1209720613;
assign addr[65164]= 1145766716;
assign addr[65165]= 1080359326;
assign addr[65166]= 1013581418;
assign addr[65167]= 945517704;
assign addr[65168]= 876254528;
assign addr[65169]= 805879757;
assign addr[65170]= 734482665;
assign addr[65171]= 662153826;
assign addr[65172]= 588984994;
assign addr[65173]= 515068990;
assign addr[65174]= 440499581;
assign addr[65175]= 365371365;
assign addr[65176]= 289779648;
assign addr[65177]= 213820322;
assign addr[65178]= 137589750;
assign addr[65179]= 61184634;
assign addr[65180]= -15298099;
assign addr[65181]= -91761426;
assign addr[65182]= -168108346;
assign addr[65183]= -244242007;
assign addr[65184]= -320065829;
assign addr[65185]= -395483624;
assign addr[65186]= -470399716;
assign addr[65187]= -544719071;
assign addr[65188]= -618347408;
assign addr[65189]= -691191324;
assign addr[65190]= -763158411;
assign addr[65191]= -834157373;
assign addr[65192]= -904098143;
assign addr[65193]= -972891995;
assign addr[65194]= -1040451659;
assign addr[65195]= -1106691431;
assign addr[65196]= -1171527280;
assign addr[65197]= -1234876957;
assign addr[65198]= -1296660098;
assign addr[65199]= -1356798326;
assign addr[65200]= -1415215352;
assign addr[65201]= -1471837070;
assign addr[65202]= -1526591649;
assign addr[65203]= -1579409630;
assign addr[65204]= -1630224009;
assign addr[65205]= -1678970324;
assign addr[65206]= -1725586737;
assign addr[65207]= -1770014111;
assign addr[65208]= -1812196087;
assign addr[65209]= -1852079154;
assign addr[65210]= -1889612716;
assign addr[65211]= -1924749160;
assign addr[65212]= -1957443913;
assign addr[65213]= -1987655498;
assign addr[65214]= -2015345591;
assign addr[65215]= -2040479063;
assign addr[65216]= -2063024031;
assign addr[65217]= -2082951896;
assign addr[65218]= -2100237377;
assign addr[65219]= -2114858546;
assign addr[65220]= -2126796855;
assign addr[65221]= -2136037160;
assign addr[65222]= -2142567738;
assign addr[65223]= -2146380306;
assign addr[65224]= -2147470025;
assign addr[65225]= -2145835515;
assign addr[65226]= -2141478848;
assign addr[65227]= -2134405552;
assign addr[65228]= -2124624598;
assign addr[65229]= -2112148396;
assign addr[65230]= -2096992772;
assign addr[65231]= -2079176953;
assign addr[65232]= -2058723538;
assign addr[65233]= -2035658475;
assign addr[65234]= -2010011024;
assign addr[65235]= -1981813720;
assign addr[65236]= -1951102334;
assign addr[65237]= -1917915825;
assign addr[65238]= -1882296293;
assign addr[65239]= -1844288924;
assign addr[65240]= -1803941934;
assign addr[65241]= -1761306505;
assign addr[65242]= -1716436725;
assign addr[65243]= -1669389513;
assign addr[65244]= -1620224553;
assign addr[65245]= -1569004214;
assign addr[65246]= -1515793473;
assign addr[65247]= -1460659832;
assign addr[65248]= -1403673233;
assign addr[65249]= -1344905966;
assign addr[65250]= -1284432584;
assign addr[65251]= -1222329801;
assign addr[65252]= -1158676398;
assign addr[65253]= -1093553126;
assign addr[65254]= -1027042599;
assign addr[65255]= -959229189;
assign addr[65256]= -890198924;
assign addr[65257]= -820039373;
assign addr[65258]= -748839539;
assign addr[65259]= -676689746;
assign addr[65260]= -603681519;
assign addr[65261]= -529907477;
assign addr[65262]= -455461206;
assign addr[65263]= -380437148;
assign addr[65264]= -304930476;
assign addr[65265]= -229036977;
assign addr[65266]= -152852926;
assign addr[65267]= -76474970;
assign addr[65268]= 0;
assign addr[65269]= 76474970;
assign addr[65270]= 152852926;
assign addr[65271]= 229036977;
assign addr[65272]= 304930476;
assign addr[65273]= 380437148;
assign addr[65274]= 455461206;
assign addr[65275]= 529907477;
assign addr[65276]= 603681519;
assign addr[65277]= 676689746;
assign addr[65278]= 748839539;
assign addr[65279]= 820039373;
assign addr[65280]= 890198924;
assign addr[65281]= 959229189;
assign addr[65282]= 1027042599;
assign addr[65283]= 1093553126;
assign addr[65284]= 1158676398;
assign addr[65285]= 1222329801;
assign addr[65286]= 1284432584;
assign addr[65287]= 1344905966;
assign addr[65288]= 1403673233;
assign addr[65289]= 1460659832;
assign addr[65290]= 1515793473;
assign addr[65291]= 1569004214;
assign addr[65292]= 1620224553;
assign addr[65293]= 1669389513;
assign addr[65294]= 1716436725;
assign addr[65295]= 1761306505;
assign addr[65296]= 1803941934;
assign addr[65297]= 1844288924;
assign addr[65298]= 1882296293;
assign addr[65299]= 1917915825;
assign addr[65300]= 1951102334;
assign addr[65301]= 1981813720;
assign addr[65302]= 2010011024;
assign addr[65303]= 2035658475;
assign addr[65304]= 2058723538;
assign addr[65305]= 2079176953;
assign addr[65306]= 2096992772;
assign addr[65307]= 2112148396;
assign addr[65308]= 2124624598;
assign addr[65309]= 2134405552;
assign addr[65310]= 2141478848;
assign addr[65311]= 2145835515;
assign addr[65312]= 2147470025;
assign addr[65313]= 2146380306;
assign addr[65314]= 2142567738;
assign addr[65315]= 2136037160;
assign addr[65316]= 2126796855;
assign addr[65317]= 2114858546;
assign addr[65318]= 2100237377;
assign addr[65319]= 2082951896;
assign addr[65320]= 2063024031;
assign addr[65321]= 2040479063;
assign addr[65322]= 2015345591;
assign addr[65323]= 1987655498;
assign addr[65324]= 1957443913;
assign addr[65325]= 1924749160;
assign addr[65326]= 1889612716;
assign addr[65327]= 1852079154;
assign addr[65328]= 1812196087;
assign addr[65329]= 1770014111;
assign addr[65330]= 1725586737;
assign addr[65331]= 1678970324;
assign addr[65332]= 1630224009;
assign addr[65333]= 1579409630;
assign addr[65334]= 1526591649;
assign addr[65335]= 1471837070;
assign addr[65336]= 1415215352;
assign addr[65337]= 1356798326;
assign addr[65338]= 1296660098;
assign addr[65339]= 1234876957;
assign addr[65340]= 1171527280;
assign addr[65341]= 1106691431;
assign addr[65342]= 1040451659;
assign addr[65343]= 972891995;
assign addr[65344]= 904098143;
assign addr[65345]= 834157373;
assign addr[65346]= 763158411;
assign addr[65347]= 691191324;
assign addr[65348]= 618347408;
assign addr[65349]= 544719071;
assign addr[65350]= 470399716;
assign addr[65351]= 395483624;
assign addr[65352]= 320065829;
assign addr[65353]= 244242007;
assign addr[65354]= 168108346;
assign addr[65355]= 91761426;
assign addr[65356]= 15298099;
assign addr[65357]= -61184634;
assign addr[65358]= -137589750;
assign addr[65359]= -213820322;
assign addr[65360]= -289779648;
assign addr[65361]= -365371365;
assign addr[65362]= -440499581;
assign addr[65363]= -515068990;
assign addr[65364]= -588984994;
assign addr[65365]= -662153826;
assign addr[65366]= -734482665;
assign addr[65367]= -805879757;
assign addr[65368]= -876254528;
assign addr[65369]= -945517704;
assign addr[65370]= -1013581418;
assign addr[65371]= -1080359326;
assign addr[65372]= -1145766716;
assign addr[65373]= -1209720613;
assign addr[65374]= -1272139887;
assign addr[65375]= -1332945355;
assign addr[65376]= -1392059879;
assign addr[65377]= -1449408469;
assign addr[65378]= -1504918373;
assign addr[65379]= -1558519173;
assign addr[65380]= -1610142873;
assign addr[65381]= -1659723983;
assign addr[65382]= -1707199606;
assign addr[65383]= -1752509516;
assign addr[65384]= -1795596234;
assign addr[65385]= -1836405100;
assign addr[65386]= -1874884346;
assign addr[65387]= -1910985158;
assign addr[65388]= -1944661739;
assign addr[65389]= -1975871368;
assign addr[65390]= -2004574453;
assign addr[65391]= -2030734582;
assign addr[65392]= -2054318569;
assign addr[65393]= -2075296495;
assign addr[65394]= -2093641749;
assign addr[65395]= -2109331059;
assign addr[65396]= -2122344521;
assign addr[65397]= -2132665626;
assign addr[65398]= -2140281282;
assign addr[65399]= -2145181827;
assign addr[65400]= -2147361045;
assign addr[65401]= -2146816171;
assign addr[65402]= -2143547897;
assign addr[65403]= -2137560369;
assign addr[65404]= -2128861181;
assign addr[65405]= -2117461370;
assign addr[65406]= -2103375398;
assign addr[65407]= -2086621133;
assign addr[65408]= -2067219829;
assign addr[65409]= -2045196100;
assign addr[65410]= -2020577882;
assign addr[65411]= -1993396407;
assign addr[65412]= -1963686155;
assign addr[65413]= -1931484818;
assign addr[65414]= -1896833245;
assign addr[65415]= -1859775393;
assign addr[65416]= -1820358275;
assign addr[65417]= -1778631892;
assign addr[65418]= -1734649179;
assign addr[65419]= -1688465931;
assign addr[65420]= -1640140734;
assign addr[65421]= -1589734894;
assign addr[65422]= -1537312353;
assign addr[65423]= -1482939614;
assign addr[65424]= -1426685652;
assign addr[65425]= -1368621831;
assign addr[65426]= -1308821808;
assign addr[65427]= -1247361445;
assign addr[65428]= -1184318708;
assign addr[65429]= -1119773573;
assign addr[65430]= -1053807919;
assign addr[65431]= -986505429;
assign addr[65432]= -917951481;
assign addr[65433]= -848233042;
assign addr[65434]= -777438554;
assign addr[65435]= -705657826;
assign addr[65436]= -632981917;
assign addr[65437]= -559503022;
assign addr[65438]= -485314355;
assign addr[65439]= -410510029;
assign addr[65440]= -335184940;
assign addr[65441]= -259434643;
assign addr[65442]= -183355234;
assign addr[65443]= -107043224;
assign addr[65444]= -30595422;
assign addr[65445]= 45891193;
assign addr[65446]= 122319591;
assign addr[65447]= 198592817;
assign addr[65448]= 274614114;
assign addr[65449]= 350287041;
assign addr[65450]= 425515602;
assign addr[65451]= 500204365;
assign addr[65452]= 574258580;
assign addr[65453]= 647584304;
assign addr[65454]= 720088517;
assign addr[65455]= 791679244;
assign addr[65456]= 862265664;
assign addr[65457]= 931758235;
assign addr[65458]= 1000068799;
assign addr[65459]= 1067110699;
assign addr[65460]= 1132798888;
assign addr[65461]= 1197050035;
assign addr[65462]= 1259782632;
assign addr[65463]= 1320917099;
assign addr[65464]= 1380375881;
assign addr[65465]= 1438083551;
assign addr[65466]= 1493966902;
assign addr[65467]= 1547955041;
assign addr[65468]= 1599979481;
assign addr[65469]= 1649974225;
assign addr[65470]= 1697875851;
assign addr[65471]= 1743623590;
assign addr[65472]= 1787159411;
assign addr[65473]= 1828428082;
assign addr[65474]= 1867377253;
assign addr[65475]= 1903957513;
assign addr[65476]= 1938122457;
assign addr[65477]= 1969828744;
assign addr[65478]= 1999036154;
assign addr[65479]= 2025707632;
assign addr[65480]= 2049809346;
assign addr[65481]= 2071310720;
assign addr[65482]= 2090184478;
assign addr[65483]= 2106406677;
assign addr[65484]= 2119956737;
assign addr[65485]= 2130817471;
assign addr[65486]= 2138975100;
assign addr[65487]= 2144419275;
assign addr[65488]= 2147143090;
assign addr[65489]= 2147143090;
assign addr[65490]= 2144419275;
assign addr[65491]= 2138975100;
assign addr[65492]= 2130817471;
assign addr[65493]= 2119956737;
assign addr[65494]= 2106406677;
assign addr[65495]= 2090184478;
assign addr[65496]= 2071310720;
assign addr[65497]= 2049809346;
assign addr[65498]= 2025707632;
assign addr[65499]= 1999036154;
assign addr[65500]= 1969828744;
assign addr[65501]= 1938122457;
assign addr[65502]= 1903957513;
assign addr[65503]= 1867377253;
assign addr[65504]= 1828428082;
assign addr[65505]= 1787159411;
assign addr[65506]= 1743623590;
assign addr[65507]= 1697875851;
assign addr[65508]= 1649974225;
assign addr[65509]= 1599979481;
assign addr[65510]= 1547955041;
assign addr[65511]= 1493966902;
assign addr[65512]= 1438083551;
assign addr[65513]= 1380375881;
assign addr[65514]= 1320917099;
assign addr[65515]= 1259782632;
assign addr[65516]= 1197050035;
assign addr[65517]= 1132798888;
assign addr[65518]= 1067110699;
assign addr[65519]= 1000068799;
assign addr[65520]= 931758235;
assign addr[65521]= 862265664;
assign addr[65522]= 791679244;
assign addr[65523]= 720088517;
assign addr[65524]= 647584304;
assign addr[65525]= 574258580;
assign addr[65526]= 500204365;
assign addr[65527]= 425515602;
assign addr[65528]= 350287041;
assign addr[65529]= 274614114;
assign addr[65530]= 198592817;
assign addr[65531]= 122319591;
assign addr[65532]= 45891193;
assign addr[65533]= -30595422;
assign addr[65534]= -107043224;
assign addr[65535]= -183355234;
endmodule